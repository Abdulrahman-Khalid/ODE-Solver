/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 21:20:01 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1415169979 */

module flipflop__2_64(D, load, Clk, Q, rst);
   input D;
   input load;
   input Clk;
   output Q;
   input rst;

   DFFR_X1 Q_reg (.D(n_0), .RN(D), .CK(n_1), .Q(Q), .QN());
   MUX2_X1 Q_reg_enable_mux_0 (.A(Q), .B(D), .S(load), .Z(n_0));
   INV_X1 i_0_0 (.A(Clk), .ZN(n_1));
endmodule

module flipflop(D, load, Clk, Q, rst);
   input D;
   input load;
   input Clk;
   output Q;
   input rst;

   DFFR_X1 Q_reg (.D(n_0), .RN(n_2), .CK(n_1), .Q(Q), .QN());
   MUX2_X1 Q_reg_enable_mux_0 (.A(Q), .B(D), .S(load), .Z(n_0));
   INV_X1 i_0_0 (.A(Clk), .ZN(n_1));
   INV_X1 i_1_0 (.A(rst), .ZN(n_2));
endmodule

module Partial_Full_Adder__2_4(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   INV_X1 i_3 (.A(P), .ZN(S));
   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_8(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_12(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_16(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_20(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_24(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_28(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_32(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_36(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_40(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_44(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_48(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_52(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_56(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_60(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_0(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire G;
   wire P;
   wire c15;
   wire n_0_0;
   wire c14;
   wire n_0_1;
   wire c13;
   wire n_0_2;
   wire c12;
   wire n_0_3;
   wire c11;
   wire n_0_4;
   wire c10;
   wire n_0_5;
   wire c9;
   wire n_0_6;
   wire c8;
   wire n_0_7;
   wire c7;
   wire n_0_8;
   wire c6;
   wire n_0_9;
   wire c5;
   wire n_0_10;
   wire c4;
   wire n_0_11;
   wire c3;
   wire n_0_12;
   wire c2;
   wire n_0_13;
   wire c1;

   Partial_Full_Adder__2_4 PFA1 (.A(A[0]), .B(B[0]), .Cin(), .S(S[0]), .P(P), 
      .G(G));
   Partial_Full_Adder__2_8 PFA2 (.A(A[1]), .B(B[1]), .Cin(c1), .S(S[1]), 
      .P(n_1), .G(n_0));
   Partial_Full_Adder__2_12 PFA3 (.A(A[2]), .B(B[2]), .Cin(c2), .S(S[2]), 
      .P(n_3), .G(n_2));
   Partial_Full_Adder__2_16 PFA4 (.A(A[3]), .B(B[3]), .Cin(c3), .S(S[3]), 
      .P(n_5), .G(n_4));
   Partial_Full_Adder__2_20 PFA5 (.A(A[4]), .B(B[4]), .Cin(c4), .S(S[4]), 
      .P(n_7), .G(n_6));
   Partial_Full_Adder__2_24 PFA6 (.A(A[5]), .B(B[5]), .Cin(c5), .S(S[5]), 
      .P(n_9), .G(n_8));
   Partial_Full_Adder__2_28 PFA7 (.A(A[6]), .B(B[6]), .Cin(c6), .S(S[6]), 
      .P(n_11), .G(n_10));
   Partial_Full_Adder__2_32 PFA8 (.A(A[7]), .B(B[7]), .Cin(c7), .S(S[7]), 
      .P(n_13), .G(n_12));
   Partial_Full_Adder__2_36 PFA9 (.A(A[8]), .B(B[8]), .Cin(c8), .S(S[8]), 
      .P(n_15), .G(n_14));
   Partial_Full_Adder__2_40 PFA10 (.A(A[9]), .B(B[9]), .Cin(c9), .S(S[9]), 
      .P(n_17), .G(n_16));
   Partial_Full_Adder__2_44 PFA11 (.A(A[10]), .B(B[10]), .Cin(c10), .S(S[10]), 
      .P(n_19), .G(n_18));
   Partial_Full_Adder__2_48 PFA12 (.A(A[11]), .B(B[11]), .Cin(c11), .S(S[11]), 
      .P(n_21), .G(n_20));
   Partial_Full_Adder__2_52 PFA13 (.A(A[12]), .B(B[12]), .Cin(c12), .S(S[12]), 
      .P(n_23), .G(n_22));
   Partial_Full_Adder__2_56 PFA14 (.A(A[13]), .B(B[13]), .Cin(c13), .S(S[13]), 
      .P(n_25), .G(n_24));
   Partial_Full_Adder__2_60 PFA15 (.A(A[14]), .B(B[14]), .Cin(c14), .S(S[14]), 
      .P(n_27), .G(n_26));
   Partial_Full_Adder__2_0 PFA16 (.A(A[15]), .B(B[15]), .Cin(c15), .S(S[15]), 
      .P(), .G());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(c15));
   AOI21_X1 i_0_1 (.A(n_26), .B1(n_27), .B2(c14), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(c14));
   AOI21_X1 i_0_3 (.A(n_24), .B1(n_25), .B2(c13), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(c13));
   AOI21_X1 i_0_5 (.A(n_22), .B1(n_23), .B2(c12), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(c12));
   AOI21_X1 i_0_7 (.A(n_20), .B1(n_21), .B2(c11), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(c11));
   AOI21_X1 i_0_9 (.A(n_18), .B1(n_19), .B2(c10), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(c10));
   AOI21_X1 i_0_11 (.A(n_16), .B1(n_17), .B2(c9), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(c9));
   AOI21_X1 i_0_13 (.A(n_14), .B1(n_15), .B2(c8), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(c8));
   AOI21_X1 i_0_15 (.A(n_12), .B1(n_13), .B2(c7), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(c7));
   AOI21_X1 i_0_17 (.A(n_10), .B1(n_11), .B2(c6), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(c6));
   AOI21_X1 i_0_19 (.A(n_8), .B1(n_9), .B2(c5), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(c5));
   AOI21_X1 i_0_21 (.A(n_6), .B1(n_7), .B2(c4), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(c4));
   AOI21_X1 i_0_23 (.A(n_4), .B1(n_5), .B2(c3), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(c3));
   AOI21_X1 i_0_25 (.A(n_2), .B1(n_3), .B2(c2), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(c2));
   AOI21_X1 i_0_27 (.A(n_0), .B1(n_1), .B2(c1), .ZN(n_0_13));
   OR2_X1 i_0_28 (.A1(P), .A2(G), .ZN(c1));
endmodule

module datapath__0_144(Index, p_0);
   input [31:0]Index;
   output [31:0]p_0;

   INV_X1 i_0 (.A(Index[0]), .ZN(p_0[0]));
   XNOR2_X1 i_1 (.A(Index[1]), .B(Index[0]), .ZN(p_0[1]));
   OR2_X1 i_2 (.A1(Index[1]), .A2(Index[0]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(Index[2]), .B(n_0), .ZN(p_0[2]));
   OR2_X1 i_4 (.A1(Index[2]), .A2(n_0), .ZN(n_1));
   XNOR2_X1 i_5 (.A(Index[3]), .B(n_1), .ZN(p_0[3]));
   OR2_X1 i_6 (.A1(Index[3]), .A2(n_1), .ZN(n_2));
   XNOR2_X1 i_7 (.A(Index[4]), .B(n_2), .ZN(p_0[4]));
   OR2_X1 i_8 (.A1(Index[4]), .A2(n_2), .ZN(n_3));
   XNOR2_X1 i_9 (.A(Index[5]), .B(n_3), .ZN(p_0[5]));
   OR2_X1 i_10 (.A1(Index[5]), .A2(n_3), .ZN(n_4));
   XNOR2_X1 i_11 (.A(Index[6]), .B(n_4), .ZN(p_0[6]));
   OR2_X1 i_12 (.A1(Index[6]), .A2(n_4), .ZN(n_5));
   XNOR2_X1 i_13 (.A(Index[7]), .B(n_5), .ZN(p_0[7]));
   OR2_X1 i_14 (.A1(Index[7]), .A2(n_5), .ZN(n_6));
   XNOR2_X1 i_15 (.A(Index[8]), .B(n_6), .ZN(p_0[8]));
   OR2_X1 i_16 (.A1(Index[8]), .A2(n_6), .ZN(n_7));
   XNOR2_X1 i_17 (.A(Index[9]), .B(n_7), .ZN(p_0[9]));
   OR2_X1 i_18 (.A1(Index[9]), .A2(n_7), .ZN(n_8));
   XNOR2_X1 i_19 (.A(Index[10]), .B(n_8), .ZN(p_0[10]));
   OR2_X1 i_20 (.A1(Index[10]), .A2(n_8), .ZN(n_9));
   XNOR2_X1 i_21 (.A(Index[11]), .B(n_9), .ZN(p_0[11]));
   OR2_X1 i_22 (.A1(Index[11]), .A2(n_9), .ZN(n_10));
   XNOR2_X1 i_23 (.A(Index[12]), .B(n_10), .ZN(p_0[12]));
   OR2_X1 i_24 (.A1(Index[12]), .A2(n_10), .ZN(n_11));
   XNOR2_X1 i_25 (.A(Index[13]), .B(n_11), .ZN(p_0[13]));
   OR2_X1 i_26 (.A1(Index[13]), .A2(n_11), .ZN(n_12));
   XNOR2_X1 i_27 (.A(Index[14]), .B(n_12), .ZN(p_0[14]));
   OR2_X1 i_28 (.A1(Index[14]), .A2(n_12), .ZN(n_13));
   XNOR2_X1 i_29 (.A(Index[15]), .B(n_13), .ZN(p_0[15]));
   OR2_X1 i_30 (.A1(Index[15]), .A2(n_13), .ZN(n_14));
   XNOR2_X1 i_31 (.A(Index[16]), .B(n_14), .ZN(p_0[16]));
   OR2_X1 i_32 (.A1(Index[16]), .A2(n_14), .ZN(n_15));
   XNOR2_X1 i_33 (.A(Index[17]), .B(n_15), .ZN(p_0[17]));
   OR2_X1 i_34 (.A1(Index[17]), .A2(n_15), .ZN(n_16));
   XNOR2_X1 i_35 (.A(Index[18]), .B(n_16), .ZN(p_0[18]));
   OR2_X1 i_36 (.A1(Index[18]), .A2(n_16), .ZN(n_17));
   XNOR2_X1 i_37 (.A(Index[19]), .B(n_17), .ZN(p_0[19]));
   OR2_X1 i_38 (.A1(Index[19]), .A2(n_17), .ZN(n_18));
   XNOR2_X1 i_39 (.A(Index[20]), .B(n_18), .ZN(p_0[20]));
   OR2_X1 i_40 (.A1(Index[20]), .A2(n_18), .ZN(n_19));
   XNOR2_X1 i_41 (.A(Index[21]), .B(n_19), .ZN(p_0[21]));
   OR2_X1 i_42 (.A1(Index[21]), .A2(n_19), .ZN(n_20));
   XNOR2_X1 i_43 (.A(Index[22]), .B(n_20), .ZN(p_0[22]));
   OR2_X1 i_44 (.A1(Index[22]), .A2(n_20), .ZN(n_21));
   XNOR2_X1 i_45 (.A(Index[23]), .B(n_21), .ZN(p_0[23]));
   OR2_X1 i_46 (.A1(Index[23]), .A2(n_21), .ZN(n_22));
   XNOR2_X1 i_47 (.A(Index[24]), .B(n_22), .ZN(p_0[24]));
   OR2_X1 i_48 (.A1(Index[24]), .A2(n_22), .ZN(n_23));
   XNOR2_X1 i_49 (.A(Index[25]), .B(n_23), .ZN(p_0[25]));
   OR2_X1 i_50 (.A1(Index[25]), .A2(n_23), .ZN(n_24));
   XNOR2_X1 i_51 (.A(Index[26]), .B(n_24), .ZN(p_0[26]));
   OR2_X1 i_52 (.A1(Index[26]), .A2(n_24), .ZN(n_25));
   XNOR2_X1 i_53 (.A(Index[27]), .B(n_25), .ZN(p_0[27]));
   OR2_X1 i_54 (.A1(Index[27]), .A2(n_25), .ZN(n_26));
   XNOR2_X1 i_55 (.A(Index[28]), .B(n_26), .ZN(p_0[28]));
   OR2_X1 i_56 (.A1(Index[28]), .A2(n_26), .ZN(n_27));
   XNOR2_X1 i_57 (.A(Index[29]), .B(n_27), .ZN(p_0[29]));
   OR2_X1 i_58 (.A1(Index[29]), .A2(n_27), .ZN(n_28));
   XNOR2_X1 i_59 (.A(Index[30]), .B(n_28), .ZN(p_0[30]));
   OR2_X1 i_60 (.A1(Index[30]), .A2(n_28), .ZN(n_29));
   XNOR2_X1 i_61 (.A(Index[31]), .B(n_29), .ZN(p_0[31]));
endmodule

module fixed_division(Dividend, Divisor, Reset, clk, Start, Quotient, ERR, Done, 
      OverFlow);
   input [15:0]Dividend;
   input [15:0]Divisor;
   input Reset;
   input clk;
   input Start;
   output [15:0]Quotient;
   output ERR;
   output Done;
   output OverFlow;

   wire [15:0]addOut;
   wire [15:0]add2;
   wire [15:0]add1;
   wire n_0_19__0;
   wire n_0_20;
   wire n_0_0;
   wire n_0_1;
   wire n_0_16;
   wire n_0_2;
   wire n_0_14__0;
   wire n_0_3;
   wire n_0_15;
   wire n_0_4__0;
   wire n_0_13;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9__0;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_17;
   wire n_0_18;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24__0;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29__0;
   wire n_0_30;
   wire n_0_31;
   wire [15:0]Dividend2;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34__0;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39__0;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44__0;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49__0;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54__0;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59__0;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64__0;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69__0;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74__0;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire [15:0]QuotientVar;
   wire [31:0]Index;
   wire n_0_123;
   wire FIRST_ONE;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_4__1;
   wire n_0_9__1;
   wire n_0_14__1;
   wire n_0_19__1;
   wire n_0_24__1;
   wire n_0_29__1;
   wire n_0_34__1;
   wire n_0_39__1;
   wire n_0_44__1;
   wire n_0_49__1;
   wire n_0_54__1;
   wire n_0_59__1;
   wire n_0_64__1;
   wire n_0_69__1;
   wire n_0_74__1;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;

   Carry_Look_Ahead u1 (.A(add1), .B(add2), .Cin(), .S(addOut));
   DLH_X1 Done_reg (.D(n_196), .G(n_194), .Q(Done));
   DLH_X1 \Quotient_reg[15]  (.D(n_193), .G(n_177), .Q(Quotient[15]));
   DLH_X1 \Quotient_reg[14]  (.D(n_192), .G(n_177), .Q(Quotient[14]));
   DLH_X1 \Quotient_reg[13]  (.D(n_191), .G(n_177), .Q(Quotient[13]));
   DLH_X1 \Quotient_reg[12]  (.D(n_190), .G(n_177), .Q(Quotient[12]));
   DLH_X1 \Quotient_reg[11]  (.D(n_189), .G(n_177), .Q(Quotient[11]));
   DLH_X1 \Quotient_reg[10]  (.D(n_188), .G(n_177), .Q(Quotient[10]));
   DLH_X1 \Quotient_reg[9]  (.D(n_187), .G(n_177), .Q(Quotient[9]));
   DLH_X1 \Quotient_reg[8]  (.D(n_186), .G(n_177), .Q(Quotient[8]));
   DLH_X1 \Quotient_reg[7]  (.D(n_185), .G(n_177), .Q(Quotient[7]));
   DLH_X1 \Quotient_reg[6]  (.D(n_184), .G(n_177), .Q(Quotient[6]));
   DLH_X1 \Quotient_reg[5]  (.D(n_183), .G(n_177), .Q(Quotient[5]));
   DLH_X1 \Quotient_reg[4]  (.D(n_182), .G(n_177), .Q(Quotient[4]));
   DLH_X1 \Quotient_reg[3]  (.D(n_181), .G(n_177), .Q(Quotient[3]));
   DLH_X1 \Quotient_reg[2]  (.D(n_180), .G(n_177), .Q(Quotient[2]));
   DLH_X1 \Quotient_reg[1]  (.D(n_179), .G(n_177), .Q(Quotient[1]));
   DLH_X1 \Quotient_reg[0]  (.D(n_178), .G(n_177), .Q(Quotient[0]));
   DLH_X1 \add2_reg[15]  (.D(n_0_74__1), .G(n_176), .Q(add2[15]));
   DLH_X1 \add2_reg[14]  (.D(n_0_69__1), .G(n_176), .Q(add2[14]));
   DLH_X1 \add2_reg[13]  (.D(n_0_64__1), .G(n_176), .Q(add2[13]));
   DLH_X1 \add2_reg[12]  (.D(n_0_59__1), .G(n_176), .Q(add2[12]));
   DLH_X1 \add2_reg[11]  (.D(n_0_54__1), .G(n_176), .Q(add2[11]));
   DLH_X1 \add2_reg[10]  (.D(n_0_49__1), .G(n_176), .Q(add2[10]));
   DLH_X1 \add2_reg[9]  (.D(n_0_44__1), .G(n_176), .Q(add2[9]));
   DLH_X1 \add2_reg[8]  (.D(n_0_39__1), .G(n_176), .Q(add2[8]));
   DLH_X1 \add2_reg[7]  (.D(n_0_34__1), .G(n_176), .Q(add2[7]));
   DLH_X1 \add2_reg[6]  (.D(n_0_29__1), .G(n_176), .Q(add2[6]));
   DLH_X1 \add2_reg[5]  (.D(n_0_24__1), .G(n_176), .Q(add2[5]));
   DLH_X1 \add2_reg[4]  (.D(n_0_19__1), .G(n_176), .Q(add2[4]));
   DLH_X1 \add2_reg[3]  (.D(n_0_14__1), .G(n_176), .Q(add2[3]));
   DLH_X1 \add2_reg[2]  (.D(n_0_9__1), .G(n_176), .Q(add2[2]));
   DLH_X1 \add2_reg[1]  (.D(n_0_4__1), .G(n_176), .Q(add2[1]));
   DLH_X1 \add2_reg[0]  (.D(n_213), .G(n_176), .Q(add2[0]));
   DLH_X1 \add1_reg[15]  (.D(n_212), .G(n_176), .Q(add1[15]));
   DLH_X1 \add1_reg[14]  (.D(n_211), .G(n_176), .Q(add1[14]));
   DLH_X1 \add1_reg[13]  (.D(n_210), .G(n_176), .Q(add1[13]));
   DLH_X1 \add1_reg[12]  (.D(n_209), .G(n_176), .Q(add1[12]));
   DLH_X1 \add1_reg[11]  (.D(n_208), .G(n_176), .Q(add1[11]));
   DLH_X1 \add1_reg[10]  (.D(n_207), .G(n_176), .Q(add1[10]));
   DLH_X1 \add1_reg[9]  (.D(n_206), .G(n_176), .Q(add1[9]));
   DLH_X1 \add1_reg[8]  (.D(n_205), .G(n_176), .Q(add1[8]));
   DLH_X1 \add1_reg[7]  (.D(n_204), .G(n_176), .Q(add1[7]));
   DLH_X1 \add1_reg[6]  (.D(n_203), .G(n_176), .Q(add1[6]));
   DLH_X1 \add1_reg[5]  (.D(n_202), .G(n_176), .Q(add1[5]));
   DLH_X1 \add1_reg[4]  (.D(n_201), .G(n_176), .Q(add1[4]));
   DLH_X1 \add1_reg[3]  (.D(n_200), .G(n_176), .Q(add1[3]));
   DLH_X1 \add1_reg[2]  (.D(n_199), .G(n_176), .Q(add1[2]));
   DLH_X1 \add1_reg[1]  (.D(n_198), .G(n_176), .Q(add1[1]));
   DLH_X1 \add1_reg[0]  (.D(n_197), .G(n_176), .Q(add1[0]));
   DLH_X1 Done_bit_reg (.D(n_175), .G(n_174), .Q(n_0));
   DLH_X1 \Index_reg[31]  (.D(Index[31]), .G(n_195), .Q(n_1));
   DLH_X1 \Index_reg[30]  (.D(Index[30]), .G(n_195), .Q(n_2));
   DLH_X1 \Index_reg[29]  (.D(Index[29]), .G(n_195), .Q(n_3));
   DLH_X1 \Index_reg[28]  (.D(Index[28]), .G(n_195), .Q(n_4));
   DLH_X1 \Index_reg[27]  (.D(Index[27]), .G(n_195), .Q(n_5));
   DLH_X1 \Index_reg[26]  (.D(Index[26]), .G(n_195), .Q(n_6));
   DLH_X1 \Index_reg[25]  (.D(Index[25]), .G(n_195), .Q(n_7));
   DLH_X1 \Index_reg[24]  (.D(Index[24]), .G(n_195), .Q(n_8));
   DLH_X1 \Index_reg[23]  (.D(Index[23]), .G(n_195), .Q(n_9));
   DLH_X1 \Index_reg[22]  (.D(Index[22]), .G(n_195), .Q(n_10));
   DLH_X1 \Index_reg[21]  (.D(Index[21]), .G(n_195), .Q(n_11));
   DLH_X1 \Index_reg[20]  (.D(Index[20]), .G(n_195), .Q(n_12));
   DLH_X1 \Index_reg[19]  (.D(Index[19]), .G(n_195), .Q(n_13));
   DLH_X1 \Index_reg[18]  (.D(Index[18]), .G(n_195), .Q(n_14));
   DLH_X1 \Index_reg[17]  (.D(Index[17]), .G(n_195), .Q(n_15));
   DLH_X1 \Index_reg[16]  (.D(Index[16]), .G(n_195), .Q(n_16));
   DLH_X1 \Index_reg[15]  (.D(Index[15]), .G(n_195), .Q(n_17));
   DLH_X1 \Index_reg[14]  (.D(Index[14]), .G(n_195), .Q(n_18));
   DLH_X1 \Index_reg[13]  (.D(Index[13]), .G(n_195), .Q(n_19));
   DLH_X1 \Index_reg[12]  (.D(Index[12]), .G(n_195), .Q(n_20));
   DLH_X1 \Index_reg[11]  (.D(Index[11]), .G(n_195), .Q(n_21));
   DLH_X1 \Index_reg[10]  (.D(Index[10]), .G(n_195), .Q(n_22));
   DLH_X1 \Index_reg[9]  (.D(Index[9]), .G(n_195), .Q(n_23));
   DLH_X1 \Index_reg[8]  (.D(Index[8]), .G(n_195), .Q(n_24));
   DLH_X1 \Index_reg[7]  (.D(Index[7]), .G(n_195), .Q(n_25));
   DLH_X1 \Index_reg[6]  (.D(Index[6]), .G(n_195), .Q(n_26));
   DLH_X1 \Index_reg[5]  (.D(Index[5]), .G(n_195), .Q(n_27));
   DLH_X1 \Index_reg[4]  (.D(Index[4]), .G(n_195), .Q(n_28));
   DLH_X1 \Index_reg[3]  (.D(Index[3]), .G(n_195), .Q(n_29));
   DLH_X1 \Index_reg[2]  (.D(Index[2]), .G(n_195), .Q(n_30));
   DLH_X1 \Index_reg[1]  (.D(Index[1]), .G(n_195), .Q(n_31));
   DLH_X1 \Index_reg[0]  (.D(Index[0]), .G(n_195), .Q(n_32));
   datapath__0_144 i_29 (.Index({n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, 
      n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, 
      n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32}), 
      .p_0({n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
      n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
      n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33}));
   DLH_X1 \QuotientVar_reg[15]  (.D(QuotientVar[15]), .G(n_173), .Q(n_65));
   DLH_X1 \QuotientVar_reg[14]  (.D(QuotientVar[14]), .G(n_172), .Q(n_66));
   DLH_X1 \QuotientVar_reg[13]  (.D(QuotientVar[13]), .G(n_171), .Q(n_67));
   DLH_X1 \QuotientVar_reg[12]  (.D(QuotientVar[12]), .G(n_170), .Q(n_68));
   DLH_X1 \QuotientVar_reg[11]  (.D(QuotientVar[11]), .G(n_169), .Q(n_69));
   DLH_X1 \QuotientVar_reg[10]  (.D(QuotientVar[10]), .G(n_168), .Q(n_70));
   DLH_X1 \QuotientVar_reg[9]  (.D(QuotientVar[9]), .G(n_167), .Q(n_71));
   DLH_X1 \QuotientVar_reg[8]  (.D(QuotientVar[8]), .G(n_166), .Q(n_72));
   DLH_X1 \QuotientVar_reg[7]  (.D(QuotientVar[7]), .G(n_165), .Q(n_73));
   DLH_X1 \QuotientVar_reg[6]  (.D(QuotientVar[6]), .G(n_164), .Q(n_74));
   DLH_X1 \QuotientVar_reg[5]  (.D(QuotientVar[5]), .G(n_163), .Q(n_75));
   DLH_X1 \QuotientVar_reg[4]  (.D(QuotientVar[4]), .G(n_162), .Q(n_76));
   DLH_X1 \QuotientVar_reg[3]  (.D(QuotientVar[3]), .G(n_161), .Q(n_77));
   DLH_X1 \QuotientVar_reg[2]  (.D(QuotientVar[2]), .G(n_160), .Q(n_78));
   DLH_X1 \QuotientVar_reg[1]  (.D(QuotientVar[1]), .G(n_159), .Q(n_79));
   DLH_X1 \QuotientVar_reg[0]  (.D(QuotientVar[0]), .G(n_158), .Q(n_80));
   DLH_X1 \Divisor2_reg[28]  (.D(n_157), .G(n_195), .Q(n_81));
   DLH_X1 \Divisor2_reg[27]  (.D(n_156), .G(n_195), .Q(n_82));
   DLH_X1 \Divisor2_reg[26]  (.D(n_155), .G(n_195), .Q(n_83));
   DLH_X1 \Divisor2_reg[25]  (.D(n_154), .G(n_195), .Q(n_84));
   DLH_X1 \Divisor2_reg[24]  (.D(n_153), .G(n_195), .Q(n_85));
   DLH_X1 \Divisor2_reg[23]  (.D(n_152), .G(n_195), .Q(n_86));
   DLH_X1 \Divisor2_reg[22]  (.D(n_151), .G(n_195), .Q(n_87));
   DLH_X1 \Divisor2_reg[21]  (.D(n_150), .G(n_195), .Q(n_88));
   DLH_X1 \Divisor2_reg[20]  (.D(n_149), .G(n_195), .Q(n_89));
   DLH_X1 \Divisor2_reg[19]  (.D(n_148), .G(n_195), .Q(n_90));
   DLH_X1 \Divisor2_reg[18]  (.D(n_147), .G(n_195), .Q(n_91));
   DLH_X1 \Divisor2_reg[17]  (.D(n_146), .G(n_195), .Q(n_92));
   DLH_X1 \Divisor2_reg[16]  (.D(n_145), .G(n_195), .Q(n_93));
   DLH_X1 \Divisor2_reg[15]  (.D(n_144), .G(n_195), .Q(n_94));
   DLH_X1 \Divisor2_reg[14]  (.D(n_143), .G(n_195), .Q(n_95));
   DLH_X1 \Divisor2_reg[13]  (.D(n_142), .G(n_195), .Q(n_96));
   DLH_X1 \Divisor2_reg[12]  (.D(n_141), .G(n_195), .Q(n_97));
   DLH_X1 \Divisor2_reg[11]  (.D(n_140), .G(n_195), .Q(n_98));
   DLH_X1 \Divisor2_reg[10]  (.D(n_139), .G(n_195), .Q(n_99));
   DLH_X1 \Divisor2_reg[9]  (.D(n_138), .G(n_195), .Q(n_100));
   DLH_X1 \Divisor2_reg[8]  (.D(n_137), .G(n_195), .Q(n_101));
   DLH_X1 \Divisor2_reg[7]  (.D(n_136), .G(n_195), .Q(n_102));
   DLH_X1 \Divisor2_reg[6]  (.D(n_135), .G(n_195), .Q(n_103));
   DLH_X1 \Divisor2_reg[5]  (.D(n_134), .G(n_195), .Q(n_104));
   DLH_X1 \Divisor2_reg[4]  (.D(n_133), .G(n_195), .Q(n_105));
   DLH_X1 \Divisor2_reg[3]  (.D(n_132), .G(n_195), .Q(n_106));
   DLH_X1 \Divisor2_reg[2]  (.D(n_131), .G(n_195), .Q(n_107));
   DLH_X1 \Divisor2_reg[1]  (.D(n_130), .G(n_195), .Q(n_108));
   DLH_X1 \Divisor2_reg[0]  (.D(n_129), .G(n_195), .Q(n_109));
   DLH_X1 \Dividend2_reg[15]  (.D(Dividend2[15]), .G(n_128), .Q(n_110));
   DLH_X1 \Dividend2_reg[14]  (.D(Dividend2[14]), .G(n_128), .Q(n_111));
   DLH_X1 \Dividend2_reg[13]  (.D(Dividend2[13]), .G(n_128), .Q(n_112));
   DLH_X1 \Dividend2_reg[12]  (.D(Dividend2[12]), .G(n_128), .Q(n_113));
   DLH_X1 \Dividend2_reg[11]  (.D(Dividend2[11]), .G(n_128), .Q(n_114));
   DLH_X1 \Dividend2_reg[10]  (.D(Dividend2[10]), .G(n_128), .Q(n_115));
   DLH_X1 \Dividend2_reg[9]  (.D(Dividend2[9]), .G(n_128), .Q(n_116));
   DLH_X1 \Dividend2_reg[8]  (.D(Dividend2[8]), .G(n_128), .Q(n_117));
   DLH_X1 \Dividend2_reg[7]  (.D(Dividend2[7]), .G(n_128), .Q(n_118));
   DLH_X1 \Dividend2_reg[6]  (.D(Dividend2[6]), .G(n_128), .Q(n_119));
   DLH_X1 \Dividend2_reg[5]  (.D(Dividend2[5]), .G(n_128), .Q(n_120));
   DLH_X1 \Dividend2_reg[4]  (.D(Dividend2[4]), .G(n_128), .Q(n_121));
   DLH_X1 \Dividend2_reg[3]  (.D(Dividend2[3]), .G(n_128), .Q(n_122));
   DLH_X1 \Dividend2_reg[2]  (.D(Dividend2[2]), .G(n_128), .Q(n_123));
   DLH_X1 \Dividend2_reg[1]  (.D(Dividend2[1]), .G(n_128), .Q(n_124));
   DLH_X1 \Dividend2_reg[0]  (.D(Dividend2[0]), .G(n_128), .Q(n_125));
   DLH_X1 FIRST_ONE_reg (.D(FIRST_ONE), .G(n_127), .Q(n_126));
   HA_X1 i_0_0 (.A(n_0_13), .B(n_0_14__0), .CO(n_0_19__0), .S());
   FA_X1 i_0_1 (.A(n_0_15), .B(n_0_16), .CI(n_0_19__0), .CO(n_0_20), .S());
   HA_X1 i_0_2 (.A(n_0_26), .B(n_0_10), .CO(n_0_0), .S());
   HA_X1 i_0_3 (.A(n_0_7), .B(n_0_0), .CO(n_0_1), .S());
   NAND2_X1 i_0_4 (.A1(n_0_2), .A2(n_0_245), .ZN(n_0_16));
   XNOR2_X1 i_0_5 (.A(n_0_253), .B(n_0_110), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(n_0_15), .A2(n_0_3), .ZN(n_0_14__0));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4__0), .ZN(n_0_3));
   OR2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4__0), .ZN(n_0_15));
   XNOR2_X1 i_0_9 (.A(n_0_253), .B(n_0_245), .ZN(n_0_4__0));
   NAND4_X1 i_0_10 (.A1(n_0_25), .A2(n_0_9__0), .A3(n_0_6), .A4(n_0_5), .ZN(
      n_0_13));
   OR2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_225), .ZN(n_0_5));
   NAND2_X1 i_0_12 (.A1(n_0_7), .A2(n_0_225), .ZN(n_0_6));
   OR3_X1 i_0_13 (.A1(Divisor[14]), .A2(n_0_8), .A3(n_0_246), .ZN(n_0_7));
   AOI21_X1 i_0_14 (.A(n_0_247), .B1(n_0_112), .B2(n_0_243), .ZN(n_0_8));
   OAI211_X1 i_0_15 (.A(n_0_232), .B(n_0_10), .C1(n_0_26), .C2(n_0_228), 
      .ZN(n_0_9__0));
   OAI21_X1 i_0_16 (.A(n_0_11), .B1(n_0_12), .B2(Divisor[14]), .ZN(n_0_10));
   OAI21_X1 i_0_17 (.A(n_0_245), .B1(n_0_21), .B2(Divisor[7]), .ZN(n_0_11));
   NOR2_X1 i_0_18 (.A1(Divisor[13]), .A2(n_0_17), .ZN(n_0_12));
   NOR2_X1 i_0_19 (.A1(Divisor[12]), .A2(n_0_18), .ZN(n_0_17));
   AOI21_X1 i_0_20 (.A(Divisor[11]), .B1(n_0_290), .B2(Divisor[9]), .ZN(n_0_18));
   NOR2_X1 i_0_21 (.A1(Divisor[6]), .A2(n_0_22), .ZN(n_0_21));
   NOR2_X1 i_0_22 (.A1(Divisor[5]), .A2(n_0_23), .ZN(n_0_22));
   NOR2_X1 i_0_23 (.A1(Divisor[4]), .A2(n_0_24__0), .ZN(n_0_23));
   AOI21_X1 i_0_24 (.A(Divisor[3]), .B1(n_0_289), .B2(Divisor[1]), .ZN(n_0_24__0));
   NAND2_X1 i_0_25 (.A1(n_0_26), .A2(n_0_228), .ZN(n_0_25));
   OAI21_X1 i_0_26 (.A(n_0_27), .B1(n_0_246), .B2(n_0_249), .ZN(n_0_26));
   AOI21_X1 i_0_27 (.A(Divisor[14]), .B1(n_0_28), .B2(n_0_245), .ZN(n_0_27));
   OR3_X1 i_0_28 (.A1(Divisor[7]), .A2(Divisor[6]), .A3(n_0_29__0), .ZN(n_0_28));
   NOR3_X1 i_0_29 (.A1(Divisor[5]), .A2(Divisor[4]), .A3(n_0_244), .ZN(n_0_29__0));
   NOR3_X1 i_0_30 (.A1(Reset), .A2(n_0_203), .A3(n_0_30), .ZN(n_127));
   NOR3_X1 i_0_31 (.A1(n_0), .A2(n_126), .A3(n_0_161), .ZN(n_0_30));
   AOI21_X1 i_0_32 (.A(Reset), .B1(n_0_105), .B2(n_0_31), .ZN(n_128));
   NAND2_X1 i_0_33 (.A1(n_0_286), .A2(n_126), .ZN(n_0_31));
   OAI21_X1 i_0_34 (.A(n_0_128), .B1(n_0_278), .B2(n_0), .ZN(Dividend2[0]));
   OAI21_X1 i_0_35 (.A(n_0_34__0), .B1(n_0_32), .B2(n_0_262), .ZN(Dividend2[1]));
   XNOR2_X1 i_0_36 (.A(n_0_293), .B(n_0_33), .ZN(n_0_32));
   NAND2_X1 i_0_37 (.A1(Dividend[15]), .A2(Dividend[0]), .ZN(n_0_33));
   NAND2_X1 i_0_38 (.A1(n_0_286), .A2(addOut[1]), .ZN(n_0_34__0));
   OAI21_X1 i_0_39 (.A(n_0_36), .B1(n_0_35), .B2(n_0_262), .ZN(Dividend2[2]));
   XNOR2_X1 i_0_40 (.A(n_0_294), .B(n_0_40), .ZN(n_0_35));
   NAND2_X1 i_0_41 (.A1(n_0_286), .A2(addOut[2]), .ZN(n_0_36));
   OAI21_X1 i_0_42 (.A(n_0_37), .B1(n_0_38), .B2(n_0_262), .ZN(Dividend2[3]));
   NAND2_X1 i_0_43 (.A1(n_0_286), .A2(addOut[3]), .ZN(n_0_37));
   XNOR2_X1 i_0_44 (.A(Dividend[3]), .B(n_0_39__0), .ZN(n_0_38));
   OAI21_X1 i_0_45 (.A(n_0_40), .B1(n_0_294), .B2(n_0_307), .ZN(n_0_39__0));
   OAI21_X1 i_0_46 (.A(Dividend[15]), .B1(Dividend[1]), .B2(Dividend[0]), 
      .ZN(n_0_40));
   OAI22_X1 i_0_47 (.A1(n_0_262), .A2(n_0_41), .B1(n_0), .B2(n_0_279), .ZN(
      Dividend2[4]));
   XNOR2_X1 i_0_48 (.A(n_0_296), .B(n_0_44__0), .ZN(n_0_41));
   OAI22_X1 i_0_49 (.A1(n_0_262), .A2(n_0_42), .B1(n_0), .B2(n_0_280), .ZN(
      Dividend2[5]));
   XNOR2_X1 i_0_50 (.A(n_0_297), .B(n_0_43), .ZN(n_0_42));
   OAI21_X1 i_0_51 (.A(Dividend[15]), .B1(n_0_261), .B2(Dividend[4]), .ZN(n_0_43));
   NAND2_X1 i_0_52 (.A1(n_0_261), .A2(Dividend[15]), .ZN(n_0_44__0));
   OAI21_X1 i_0_53 (.A(n_0_46), .B1(n_0_45), .B2(n_0_262), .ZN(Dividend2[6]));
   XNOR2_X1 i_0_54 (.A(n_0_298), .B(n_0_50), .ZN(n_0_45));
   NAND2_X1 i_0_55 (.A1(n_0_286), .A2(addOut[6]), .ZN(n_0_46));
   OAI21_X1 i_0_56 (.A(n_0_48), .B1(n_0_47), .B2(n_0_262), .ZN(Dividend2[7]));
   XNOR2_X1 i_0_57 (.A(n_0_299), .B(n_0_49__0), .ZN(n_0_47));
   NAND2_X1 i_0_58 (.A1(n_0_286), .A2(addOut[7]), .ZN(n_0_48));
   OAI21_X1 i_0_59 (.A(Dividend[15]), .B1(n_0_259), .B2(Dividend[6]), .ZN(
      n_0_49__0));
   NAND2_X1 i_0_60 (.A1(n_0_259), .A2(Dividend[15]), .ZN(n_0_50));
   OAI22_X1 i_0_61 (.A1(n_0_262), .A2(n_0_51), .B1(n_0), .B2(n_0_281), .ZN(
      Dividend2[8]));
   XNOR2_X1 i_0_62 (.A(n_0_300), .B(n_0_68), .ZN(n_0_51));
   OAI22_X1 i_0_63 (.A1(n_0_262), .A2(n_0_52), .B1(n_0), .B2(n_0_282), .ZN(
      Dividend2[9]));
   XNOR2_X1 i_0_64 (.A(n_0_301), .B(n_0_53), .ZN(n_0_52));
   OAI21_X1 i_0_65 (.A(Dividend[15]), .B1(n_0_257), .B2(Dividend[8]), .ZN(n_0_53));
   OAI21_X1 i_0_66 (.A(n_0_55), .B1(n_0_54__0), .B2(n_0_262), .ZN(Dividend2[10]));
   XNOR2_X1 i_0_67 (.A(n_0_302), .B(n_0_59__0), .ZN(n_0_54__0));
   NAND2_X1 i_0_68 (.A1(n_0_286), .A2(addOut[10]), .ZN(n_0_55));
   OAI21_X1 i_0_69 (.A(n_0_57), .B1(n_0_56), .B2(n_0_262), .ZN(Dividend2[11]));
   XNOR2_X1 i_0_70 (.A(n_0_303), .B(n_0_58), .ZN(n_0_56));
   NAND2_X1 i_0_71 (.A1(n_0_286), .A2(addOut[11]), .ZN(n_0_57));
   OAI21_X1 i_0_72 (.A(Dividend[15]), .B1(n_0_252), .B2(Dividend[10]), .ZN(
      n_0_58));
   NAND2_X1 i_0_73 (.A1(n_0_252), .A2(Dividend[15]), .ZN(n_0_59__0));
   OAI22_X1 i_0_74 (.A1(n_0_262), .A2(n_0_60), .B1(n_0), .B2(n_0_283), .ZN(
      Dividend2[12]));
   XNOR2_X1 i_0_75 (.A(n_0_304), .B(n_0_67), .ZN(n_0_60));
   OAI21_X1 i_0_76 (.A(n_0_62), .B1(n_0_61), .B2(n_0_262), .ZN(Dividend2[13]));
   XNOR2_X1 i_0_77 (.A(n_0_305), .B(n_0_63), .ZN(n_0_61));
   NAND2_X1 i_0_78 (.A1(n_0_286), .A2(addOut[13]), .ZN(n_0_62));
   OAI21_X1 i_0_79 (.A(Dividend[15]), .B1(n_0_251), .B2(Dividend[12]), .ZN(
      n_0_63));
   OAI21_X1 i_0_80 (.A(n_0_65), .B1(n_0_64__0), .B2(n_0_262), .ZN(Dividend2[14]));
   XNOR2_X1 i_0_81 (.A(Dividend[14]), .B(n_0_66), .ZN(n_0_64__0));
   NAND2_X1 i_0_82 (.A1(n_0_286), .A2(addOut[14]), .ZN(n_0_65));
   OAI21_X1 i_0_83 (.A(n_0_67), .B1(n_0_256), .B2(n_0_307), .ZN(n_0_66));
   NAND2_X1 i_0_84 (.A1(n_0_251), .A2(Dividend[15]), .ZN(n_0_67));
   NAND2_X1 i_0_85 (.A1(n_0_257), .A2(Dividend[15]), .ZN(n_0_68));
   OAI21_X1 i_0_86 (.A(n_0_69__0), .B1(n_0_284), .B2(n_0), .ZN(Dividend2[15]));
   NAND3_X1 i_0_87 (.A1(Dividend[15]), .A2(n_0_313), .A3(n_0_250), .ZN(n_0_69__0));
   NOR2_X1 i_0_88 (.A1(n_0_4__1), .A2(n_0), .ZN(n_129));
   NOR2_X1 i_0_89 (.A1(n_0_9__1), .A2(n_0), .ZN(n_130));
   NOR2_X1 i_0_90 (.A1(n_0_14__1), .A2(n_0), .ZN(n_131));
   NOR2_X1 i_0_91 (.A1(n_0_19__1), .A2(n_0), .ZN(n_132));
   NOR2_X1 i_0_92 (.A1(n_0_24__1), .A2(n_0), .ZN(n_133));
   NOR2_X1 i_0_93 (.A1(n_0_29__1), .A2(n_0), .ZN(n_134));
   NOR2_X1 i_0_94 (.A1(n_0_34__1), .A2(n_0), .ZN(n_135));
   NOR2_X1 i_0_95 (.A1(n_0_39__1), .A2(n_0), .ZN(n_136));
   NOR2_X1 i_0_96 (.A1(n_0_44__1), .A2(n_0), .ZN(n_137));
   NOR2_X1 i_0_97 (.A1(n_0_49__1), .A2(n_0), .ZN(n_138));
   NOR2_X1 i_0_98 (.A1(n_0_54__1), .A2(n_0), .ZN(n_139));
   NOR2_X1 i_0_99 (.A1(n_0_59__1), .A2(n_0), .ZN(n_140));
   NOR2_X1 i_0_100 (.A1(n_0_64__1), .A2(n_0), .ZN(n_141));
   NOR2_X1 i_0_101 (.A1(n_0_69__1), .A2(n_0), .ZN(n_142));
   OAI22_X1 i_0_102 (.A1(n_0_287), .A2(n_0_105), .B1(n_0), .B2(n_0_74__1), 
      .ZN(n_143));
   OAI21_X1 i_0_103 (.A(n_0_72), .B1(n_0_105), .B2(n_0_70), .ZN(n_144));
   XNOR2_X1 i_0_104 (.A(n_0_288), .B(n_0_71), .ZN(n_0_70));
   NAND2_X1 i_0_105 (.A1(Divisor[15]), .A2(Divisor[0]), .ZN(n_0_71));
   NAND2_X1 i_0_106 (.A1(n_0_286), .A2(n_93), .ZN(n_0_72));
   OAI22_X1 i_0_107 (.A1(n_0_105), .A2(n_0_73), .B1(n_0_309), .B2(n_0), .ZN(
      n_145));
   XNOR2_X1 i_0_108 (.A(n_0_289), .B(n_0_76), .ZN(n_0_73));
   OAI22_X1 i_0_109 (.A1(n_0_105), .A2(n_0_74__0), .B1(n_0_310), .B2(n_0), 
      .ZN(n_146));
   XNOR2_X1 i_0_110 (.A(Divisor[3]), .B(n_0_75), .ZN(n_0_74__0));
   OAI21_X1 i_0_111 (.A(n_0_76), .B1(n_0_289), .B2(n_0_291), .ZN(n_0_75));
   OAI21_X1 i_0_112 (.A(Divisor[15]), .B1(Divisor[1]), .B2(Divisor[0]), .ZN(
      n_0_76));
   OAI21_X1 i_0_113 (.A(n_0_78), .B1(n_0_105), .B2(n_0_77), .ZN(n_147));
   XOR2_X1 i_0_114 (.A(Divisor[4]), .B(n_0_81), .Z(n_0_77));
   NAND2_X1 i_0_115 (.A1(n_0_286), .A2(n_90), .ZN(n_0_78));
   OAI22_X1 i_0_116 (.A1(n_0_105), .A2(n_0_79), .B1(n_0_311), .B2(n_0), .ZN(
      n_148));
   XOR2_X1 i_0_117 (.A(Divisor[5]), .B(n_0_80), .Z(n_0_79));
   OAI21_X1 i_0_118 (.A(Divisor[15]), .B1(n_0_243), .B2(Divisor[4]), .ZN(n_0_80));
   NAND2_X1 i_0_119 (.A1(n_0_243), .A2(Divisor[15]), .ZN(n_0_81));
   OAI22_X1 i_0_120 (.A1(n_0_105), .A2(n_0_82), .B1(n_0_312), .B2(n_0), .ZN(
      n_149));
   XOR2_X1 i_0_121 (.A(Divisor[6]), .B(n_0_83), .Z(n_0_82));
   NAND2_X1 i_0_122 (.A1(n_0_242), .A2(Divisor[15]), .ZN(n_0_83));
   OAI21_X1 i_0_123 (.A(n_0_86), .B1(n_0_84), .B2(n_0_105), .ZN(n_150));
   XOR2_X1 i_0_124 (.A(Divisor[7]), .B(n_0_85), .Z(n_0_84));
   NAND2_X1 i_0_125 (.A1(n_0_241), .A2(Divisor[15]), .ZN(n_0_85));
   NAND2_X1 i_0_126 (.A1(n_0_286), .A2(n_87), .ZN(n_0_86));
   OAI21_X1 i_0_127 (.A(n_0_88), .B1(n_0_87), .B2(n_0_105), .ZN(n_151));
   XNOR2_X1 i_0_128 (.A(Divisor[8]), .B(n_0_97), .ZN(n_0_87));
   NAND2_X1 i_0_129 (.A1(n_0_286), .A2(n_86), .ZN(n_0_88));
   OAI21_X1 i_0_130 (.A(n_0_90), .B1(n_0_89), .B2(n_0_105), .ZN(n_152));
   XOR2_X1 i_0_131 (.A(Divisor[9]), .B(n_0_96), .Z(n_0_89));
   NAND2_X1 i_0_132 (.A1(n_0_286), .A2(n_85), .ZN(n_0_90));
   OAI21_X1 i_0_133 (.A(n_0_92), .B1(n_0_91), .B2(n_0_105), .ZN(n_153));
   XNOR2_X1 i_0_134 (.A(n_0_290), .B(n_0_95), .ZN(n_0_91));
   NAND2_X1 i_0_135 (.A1(n_0_286), .A2(n_84), .ZN(n_0_92));
   OAI21_X1 i_0_136 (.A(n_0_98), .B1(n_0_93), .B2(n_0_105), .ZN(n_154));
   XOR2_X1 i_0_137 (.A(Divisor[11]), .B(n_0_94), .Z(n_0_93));
   OAI21_X1 i_0_138 (.A(Divisor[15]), .B1(n_0_109), .B2(Divisor[10]), .ZN(n_0_94));
   NAND2_X1 i_0_139 (.A1(n_0_109), .A2(Divisor[15]), .ZN(n_0_95));
   OAI21_X1 i_0_140 (.A(Divisor[15]), .B1(n_0_110), .B2(Divisor[8]), .ZN(n_0_96));
   NOR2_X1 i_0_141 (.A1(n_0_111), .A2(n_0_291), .ZN(n_0_97));
   NAND2_X1 i_0_142 (.A1(n_0_286), .A2(n_83), .ZN(n_0_98));
   OAI21_X1 i_0_143 (.A(n_0_100), .B1(n_0_99), .B2(n_0_105), .ZN(n_155));
   XOR2_X1 i_0_144 (.A(Divisor[12]), .B(n_0_107), .Z(n_0_99));
   NAND2_X1 i_0_145 (.A1(n_0_286), .A2(n_82), .ZN(n_0_100));
   OAI21_X1 i_0_146 (.A(n_0_103), .B1(n_0_101), .B2(n_0_105), .ZN(n_156));
   XOR2_X1 i_0_147 (.A(Divisor[13]), .B(n_0_102), .Z(n_0_101));
   OAI21_X1 i_0_148 (.A(Divisor[15]), .B1(n_0_108), .B2(Divisor[12]), .ZN(
      n_0_102));
   NAND2_X1 i_0_149 (.A1(n_0_286), .A2(n_81), .ZN(n_0_103));
   NOR2_X1 i_0_150 (.A1(n_0_105), .A2(n_0_104), .ZN(n_157));
   XOR2_X1 i_0_151 (.A(Divisor[14]), .B(n_0_106), .Z(n_0_104));
   NAND2_X1 i_0_152 (.A1(n_0_313), .A2(n_0_239), .ZN(n_0_105));
   OAI21_X1 i_0_153 (.A(Divisor[15]), .B1(n_0_246), .B2(n_0_108), .ZN(n_0_106));
   NAND2_X1 i_0_154 (.A1(n_0_108), .A2(Divisor[15]), .ZN(n_0_107));
   NAND3_X1 i_0_155 (.A1(n_0_249), .A2(n_0_248), .A3(n_0_111), .ZN(n_0_108));
   NAND2_X1 i_0_156 (.A1(n_0_248), .A2(n_0_111), .ZN(n_0_109));
   INV_X1 i_0_157 (.A(n_0_111), .ZN(n_0_110));
   NOR2_X1 i_0_158 (.A1(n_0_241), .A2(Divisor[7]), .ZN(n_0_111));
   NOR4_X1 i_0_159 (.A1(Divisor[7]), .A2(Divisor[6]), .A3(Divisor[5]), .A4(
      Divisor[4]), .ZN(n_0_112));
   OAI21_X1 i_0_160 (.A(n_0_122), .B1(n_0_115), .B2(n_0_206), .ZN(n_158));
   OAI21_X1 i_0_161 (.A(n_0_122), .B1(n_0_116), .B2(n_0_206), .ZN(n_159));
   OAI21_X1 i_0_162 (.A(n_0_122), .B1(n_0_118), .B2(n_0_206), .ZN(n_160));
   OAI21_X1 i_0_163 (.A(n_0_122), .B1(n_0_119), .B2(n_0_206), .ZN(n_161));
   OAI21_X1 i_0_164 (.A(n_0_122), .B1(n_0_115), .B2(n_0_113), .ZN(n_162));
   OAI21_X1 i_0_165 (.A(n_0_122), .B1(n_0_116), .B2(n_0_113), .ZN(n_163));
   OAI21_X1 i_0_166 (.A(n_0_122), .B1(n_0_118), .B2(n_0_113), .ZN(n_164));
   OAI21_X1 i_0_167 (.A(n_0_122), .B1(n_0_119), .B2(n_0_113), .ZN(n_165));
   OR3_X1 i_0_168 (.A1(n_0_207), .A2(n_29), .A3(n_0_308), .ZN(n_0_113));
   OAI21_X1 i_0_169 (.A(n_0_122), .B1(n_0_115), .B2(n_0_114), .ZN(n_166));
   OAI21_X1 i_0_170 (.A(n_0_122), .B1(n_0_116), .B2(n_0_114), .ZN(n_167));
   OAI21_X1 i_0_171 (.A(n_0_122), .B1(n_0_118), .B2(n_0_114), .ZN(n_168));
   OAI21_X1 i_0_172 (.A(n_0_122), .B1(n_0_119), .B2(n_0_114), .ZN(n_169));
   NAND3_X1 i_0_173 (.A1(n_29), .A2(n_0_208), .A3(n_0_308), .ZN(n_0_114));
   OAI21_X1 i_0_174 (.A(n_0_122), .B1(n_0_121), .B2(n_0_115), .ZN(n_170));
   NAND2_X1 i_0_175 (.A1(n_33), .A2(n_0_117), .ZN(n_0_115));
   OAI21_X1 i_0_176 (.A(n_0_122), .B1(n_0_121), .B2(n_0_116), .ZN(n_171));
   NAND2_X1 i_0_177 (.A1(n_32), .A2(n_0_117), .ZN(n_0_116));
   NOR2_X1 i_0_178 (.A1(n_0_123), .A2(n_31), .ZN(n_0_117));
   OAI21_X1 i_0_179 (.A(n_0_122), .B1(n_0_121), .B2(n_0_118), .ZN(n_172));
   NAND2_X1 i_0_180 (.A1(n_33), .A2(n_0_120), .ZN(n_0_118));
   OAI21_X1 i_0_181 (.A(n_0_122), .B1(n_0_121), .B2(n_0_119), .ZN(n_173));
   NAND2_X1 i_0_182 (.A1(n_32), .A2(n_0_120), .ZN(n_0_119));
   AND2_X1 i_0_183 (.A1(n_31), .A2(n_176), .ZN(n_0_120));
   NAND3_X1 i_0_184 (.A1(n_29), .A2(n_30), .A3(n_0_208), .ZN(n_0_121));
   NAND2_X1 i_0_185 (.A1(n_0_313), .A2(n_0_285), .ZN(n_0_122));
   OAI21_X1 i_0_186 (.A(n_0), .B1(n_0_125), .B2(n_0_292), .ZN(QuotientVar[0]));
   OAI21_X1 i_0_187 (.A(n_0), .B1(n_0_125), .B2(n_0_293), .ZN(QuotientVar[1]));
   OAI21_X1 i_0_188 (.A(n_0), .B1(n_0_125), .B2(n_0_294), .ZN(QuotientVar[2]));
   OAI21_X1 i_0_189 (.A(n_0), .B1(n_0_125), .B2(n_0_295), .ZN(QuotientVar[3]));
   OAI21_X1 i_0_190 (.A(n_0), .B1(n_0_125), .B2(n_0_296), .ZN(QuotientVar[4]));
   OAI21_X1 i_0_191 (.A(n_0), .B1(n_0_125), .B2(n_0_297), .ZN(QuotientVar[5]));
   OAI21_X1 i_0_192 (.A(n_0), .B1(n_0_125), .B2(n_0_298), .ZN(QuotientVar[6]));
   OAI21_X1 i_0_193 (.A(n_0), .B1(n_0_125), .B2(n_0_299), .ZN(QuotientVar[7]));
   OAI21_X1 i_0_194 (.A(n_0), .B1(n_0_125), .B2(n_0_300), .ZN(QuotientVar[8]));
   OAI21_X1 i_0_195 (.A(n_0), .B1(n_0_125), .B2(n_0_301), .ZN(QuotientVar[9]));
   OAI21_X1 i_0_196 (.A(n_0), .B1(n_0_125), .B2(n_0_302), .ZN(QuotientVar[10]));
   OAI21_X1 i_0_197 (.A(n_0), .B1(n_0_125), .B2(n_0_303), .ZN(QuotientVar[11]));
   OAI21_X1 i_0_198 (.A(n_0), .B1(n_0_125), .B2(n_0_304), .ZN(QuotientVar[12]));
   OAI21_X1 i_0_199 (.A(n_0), .B1(n_0_125), .B2(n_0_305), .ZN(QuotientVar[13]));
   OAI21_X1 i_0_200 (.A(n_0), .B1(n_0_125), .B2(n_0_306), .ZN(QuotientVar[14]));
   OAI21_X1 i_0_201 (.A(n_0_262), .B1(n_0), .B2(n_32), .ZN(Index[0]));
   AND2_X1 i_0_202 (.A1(n_0_286), .A2(n_34), .ZN(Index[1]));
   OAI21_X1 i_0_203 (.A(n_0_262), .B1(n_0_271), .B2(n_0), .ZN(Index[2]));
   AND2_X1 i_0_204 (.A1(n_0_286), .A2(n_36), .ZN(Index[3]));
   OAI21_X1 i_0_205 (.A(n_0_262), .B1(n_0_272), .B2(n_0), .ZN(Index[4]));
   AND2_X1 i_0_206 (.A1(n_0_286), .A2(n_38), .ZN(Index[5]));
   AND2_X1 i_0_207 (.A1(n_0_286), .A2(n_39), .ZN(Index[6]));
   AND2_X1 i_0_208 (.A1(n_0_286), .A2(n_40), .ZN(Index[7]));
   AND2_X1 i_0_209 (.A1(n_0_286), .A2(n_41), .ZN(Index[8]));
   AND2_X1 i_0_210 (.A1(n_0_286), .A2(n_42), .ZN(Index[9]));
   AND2_X1 i_0_211 (.A1(n_0_286), .A2(n_43), .ZN(Index[10]));
   AND2_X1 i_0_212 (.A1(n_0_286), .A2(n_44), .ZN(Index[11]));
   AND2_X1 i_0_213 (.A1(n_0_286), .A2(n_45), .ZN(Index[12]));
   AND2_X1 i_0_214 (.A1(n_0_286), .A2(n_46), .ZN(Index[13]));
   AND2_X1 i_0_215 (.A1(n_0_286), .A2(n_47), .ZN(Index[14]));
   AND2_X1 i_0_216 (.A1(n_0_286), .A2(n_48), .ZN(Index[15]));
   AND2_X1 i_0_217 (.A1(n_0_286), .A2(n_49), .ZN(Index[16]));
   AND2_X1 i_0_218 (.A1(n_0_286), .A2(n_50), .ZN(Index[17]));
   AND2_X1 i_0_219 (.A1(n_0_286), .A2(n_51), .ZN(Index[18]));
   AND2_X1 i_0_220 (.A1(n_0_286), .A2(n_52), .ZN(Index[19]));
   AND2_X1 i_0_221 (.A1(n_0_286), .A2(n_53), .ZN(Index[20]));
   AND2_X1 i_0_222 (.A1(n_0_286), .A2(n_54), .ZN(Index[21]));
   AND2_X1 i_0_223 (.A1(n_0_286), .A2(n_55), .ZN(Index[22]));
   AND2_X1 i_0_224 (.A1(n_0_286), .A2(n_56), .ZN(Index[23]));
   AND2_X1 i_0_225 (.A1(n_0_286), .A2(n_57), .ZN(Index[24]));
   AND2_X1 i_0_226 (.A1(n_0_286), .A2(n_58), .ZN(Index[25]));
   AND2_X1 i_0_227 (.A1(n_0_286), .A2(n_59), .ZN(Index[26]));
   AND2_X1 i_0_228 (.A1(n_0_286), .A2(n_60), .ZN(Index[27]));
   AND2_X1 i_0_229 (.A1(n_0_286), .A2(n_61), .ZN(Index[28]));
   AND2_X1 i_0_230 (.A1(n_0_286), .A2(n_62), .ZN(Index[29]));
   AND2_X1 i_0_231 (.A1(n_0_286), .A2(n_63), .ZN(Index[30]));
   AND2_X1 i_0_232 (.A1(n_0_286), .A2(n_64), .ZN(Index[31]));
   NAND2_X1 i_0_233 (.A1(n_0_203), .A2(n_0_285), .ZN(n_174));
   OAI211_X1 i_0_234 (.A(n_0_285), .B(n_0_204), .C1(n_0_222), .C2(n_0_262), 
      .ZN(n_175));
   INV_X1 i_0_235 (.A(n_0_123), .ZN(n_176));
   NAND2_X1 i_0_236 (.A1(FIRST_ONE), .A2(n_0_285), .ZN(n_0_123));
   INV_X1 i_0_237 (.A(n_0_124), .ZN(FIRST_ONE));
   NAND2_X1 i_0_238 (.A1(n_0_161), .A2(n_0_286), .ZN(n_0_124));
   AOI21_X1 i_0_239 (.A(Reset), .B1(n_0_204), .B2(n_0_125), .ZN(n_177));
   OAI21_X1 i_0_240 (.A(n_0_313), .B1(n_0_250), .B2(n_0_126), .ZN(n_0_125));
   NOR3_X1 i_0_241 (.A1(n_0_241), .A2(n_0_127), .A3(Divisor[15]), .ZN(n_0_126));
   NAND2_X1 i_0_242 (.A1(Divisor[7]), .A2(n_0_245), .ZN(n_0_127));
   OAI21_X1 i_0_243 (.A(n_0_128), .B1(n_0_160), .B2(n_0), .ZN(n_178));
   NAND2_X1 i_0_244 (.A1(Dividend[0]), .A2(n_0_313), .ZN(n_0_128));
   OAI22_X1 i_0_245 (.A1(n_0_129), .A2(n_0), .B1(n_0_293), .B2(n_0_262), 
      .ZN(n_179));
   XNOR2_X1 i_0_246 (.A(n_79), .B(n_0_159), .ZN(n_0_129));
   OAI22_X1 i_0_247 (.A1(n_0_130), .A2(n_0), .B1(n_0_294), .B2(n_0_262), 
      .ZN(n_180));
   XOR2_X1 i_0_248 (.A(n_78), .B(n_0_158), .Z(n_0_130));
   OAI22_X1 i_0_249 (.A1(n_0_131), .A2(n_0), .B1(n_0_295), .B2(n_0_262), 
      .ZN(n_181));
   XOR2_X1 i_0_250 (.A(n_77), .B(n_0_156), .Z(n_0_131));
   OAI22_X1 i_0_251 (.A1(n_0_132), .A2(n_0), .B1(n_0_296), .B2(n_0_262), 
      .ZN(n_182));
   XNOR2_X1 i_0_252 (.A(n_76), .B(n_0_155), .ZN(n_0_132));
   OAI22_X1 i_0_253 (.A1(n_0_133), .A2(n_0), .B1(n_0_297), .B2(n_0_262), 
      .ZN(n_183));
   XNOR2_X1 i_0_254 (.A(n_75), .B(n_0_154), .ZN(n_0_133));
   OAI22_X1 i_0_255 (.A1(n_0_134), .A2(n_0), .B1(n_0_298), .B2(n_0_262), 
      .ZN(n_184));
   XNOR2_X1 i_0_256 (.A(n_0_274), .B(n_0_153), .ZN(n_0_134));
   OAI22_X1 i_0_257 (.A1(n_0_135), .A2(n_0), .B1(n_0_299), .B2(n_0_262), 
      .ZN(n_185));
   XNOR2_X1 i_0_258 (.A(n_73), .B(n_0_152), .ZN(n_0_135));
   OAI22_X1 i_0_259 (.A1(n_0_136), .A2(n_0), .B1(n_0_300), .B2(n_0_262), 
      .ZN(n_186));
   XNOR2_X1 i_0_260 (.A(n_72), .B(n_0_150), .ZN(n_0_136));
   OAI22_X1 i_0_261 (.A1(n_0_137), .A2(n_0), .B1(n_0_301), .B2(n_0_262), 
      .ZN(n_187));
   XNOR2_X1 i_0_262 (.A(n_0_275), .B(n_0_149), .ZN(n_0_137));
   OAI22_X1 i_0_263 (.A1(n_0_138), .A2(n_0), .B1(n_0_302), .B2(n_0_262), 
      .ZN(n_188));
   XNOR2_X1 i_0_264 (.A(n_70), .B(n_0_148), .ZN(n_0_138));
   OAI22_X1 i_0_265 (.A1(n_0_139), .A2(n_0), .B1(n_0_303), .B2(n_0_262), 
      .ZN(n_189));
   XNOR2_X1 i_0_266 (.A(n_69), .B(n_0_146), .ZN(n_0_139));
   OAI22_X1 i_0_267 (.A1(n_0_140), .A2(n_0), .B1(n_0_304), .B2(n_0_262), 
      .ZN(n_190));
   XNOR2_X1 i_0_268 (.A(n_0_276), .B(n_0_145), .ZN(n_0_140));
   OAI22_X1 i_0_269 (.A1(n_0_141), .A2(n_0), .B1(n_0_305), .B2(n_0_262), 
      .ZN(n_191));
   XNOR2_X1 i_0_270 (.A(n_67), .B(n_0_144), .ZN(n_0_141));
   OAI22_X1 i_0_271 (.A1(n_0_142), .A2(n_0), .B1(n_0_306), .B2(n_0_262), 
      .ZN(n_192));
   XOR2_X1 i_0_272 (.A(n_66), .B(n_0_143), .Z(n_0_142));
   AOI21_X1 i_0_273 (.A(n_0_144), .B1(n_0_200), .B2(n_67), .ZN(n_0_143));
   OAI21_X1 i_0_274 (.A(n_0_145), .B1(n_0_199), .B2(n_0_276), .ZN(n_0_144));
   AOI21_X1 i_0_275 (.A(n_0_146), .B1(n_0_200), .B2(n_69), .ZN(n_0_145));
   INV_X1 i_0_276 (.A(n_0_147), .ZN(n_0_146));
   AOI21_X1 i_0_277 (.A(n_0_148), .B1(n_0_200), .B2(n_70), .ZN(n_0_147));
   OAI21_X1 i_0_278 (.A(n_0_149), .B1(n_0_199), .B2(n_0_275), .ZN(n_0_148));
   AOI21_X1 i_0_279 (.A(n_0_150), .B1(n_0_200), .B2(n_72), .ZN(n_0_149));
   INV_X1 i_0_280 (.A(n_0_151), .ZN(n_0_150));
   AOI21_X1 i_0_281 (.A(n_0_152), .B1(n_0_200), .B2(n_73), .ZN(n_0_151));
   OAI21_X1 i_0_282 (.A(n_0_153), .B1(n_0_199), .B2(n_0_274), .ZN(n_0_152));
   AOI21_X1 i_0_283 (.A(n_0_154), .B1(n_0_200), .B2(n_75), .ZN(n_0_153));
   NAND3_X1 i_0_284 (.A1(n_0_198), .A2(n_0_197), .A3(n_0_156), .ZN(n_0_154));
   NAND2_X1 i_0_285 (.A1(n_0_197), .A2(n_0_156), .ZN(n_0_155));
   OAI21_X1 i_0_286 (.A(n_0_200), .B1(n_0_157), .B2(n_78), .ZN(n_0_156));
   NAND2_X1 i_0_287 (.A1(n_0_160), .A2(n_0_273), .ZN(n_0_157));
   AOI21_X1 i_0_288 (.A(n_0_159), .B1(n_0_200), .B2(n_79), .ZN(n_0_158));
   NOR2_X1 i_0_289 (.A1(n_0_160), .A2(n_0_199), .ZN(n_0_159));
   NOR2_X1 i_0_290 (.A1(n_80), .A2(n_0_161), .ZN(n_0_160));
   INV_X1 i_0_291 (.A(n_0_162), .ZN(n_0_161));
   NAND3_X1 i_0_292 (.A1(n_0_174), .A2(n_0_169), .A3(n_0_163), .ZN(n_0_162));
   AOI21_X1 i_0_293 (.A(n_0_164), .B1(n_0_269), .B2(n_94), .ZN(n_0_163));
   NAND4_X1 i_0_294 (.A1(n_0_168), .A2(n_0_167), .A3(n_0_166), .A4(n_0_165), 
      .ZN(n_0_164));
   NOR4_X1 i_0_295 (.A1(n_87), .A2(n_90), .A3(n_91), .A4(n_93), .ZN(n_0_165));
   NOR3_X1 i_0_296 (.A1(n_88), .A2(n_89), .A3(n_92), .ZN(n_0_166));
   NOR4_X1 i_0_297 (.A1(n_83), .A2(n_84), .A3(n_85), .A4(n_86), .ZN(n_0_167));
   NOR2_X1 i_0_298 (.A1(n_81), .A2(n_82), .ZN(n_0_168));
   NAND4_X1 i_0_299 (.A1(n_0_173), .A2(n_0_172), .A3(n_0_171), .A4(n_0_170), 
      .ZN(n_0_169));
   NOR4_X1 i_0_300 (.A1(n_200), .A2(n_199), .A3(n_198), .A4(n_197), .ZN(n_0_170));
   NOR4_X1 i_0_301 (.A1(n_204), .A2(n_203), .A3(n_202), .A4(n_201), .ZN(n_0_171));
   NOR4_X1 i_0_302 (.A1(n_208), .A2(n_207), .A3(n_206), .A4(n_205), .ZN(n_0_172));
   NOR4_X1 i_0_303 (.A1(n_211), .A2(n_210), .A3(n_209), .A4(n_212), .ZN(n_0_173));
   OAI21_X1 i_0_304 (.A(n_0_175), .B1(n_0_177), .B2(n_0_176), .ZN(n_0_174));
   AOI22_X1 i_0_305 (.A1(n_211), .A2(n_0_69__1), .B1(n_0_74__1), .B2(n_212), 
      .ZN(n_0_175));
   OAI22_X1 i_0_306 (.A1(n_0_69__1), .A2(n_211), .B1(n_210), .B2(n_0_64__1), 
      .ZN(n_0_176));
   AOI221_X1 i_0_307 (.A(n_0_178), .B1(n_209), .B2(n_0_59__1), .C1(n_0_64__1), 
      .C2(n_210), .ZN(n_0_177));
   AOI21_X1 i_0_308 (.A(n_0_179), .B1(n_0_181), .B2(n_0_180), .ZN(n_0_178));
   OAI22_X1 i_0_309 (.A1(n_0_54__1), .A2(n_208), .B1(n_209), .B2(n_0_59__1), 
      .ZN(n_0_179));
   AOI22_X1 i_0_310 (.A1(n_0_54__1), .A2(n_208), .B1(n_207), .B2(n_0_49__1), 
      .ZN(n_0_180));
   OR2_X1 i_0_311 (.A1(n_0_183), .A2(n_0_182), .ZN(n_0_181));
   OAI22_X1 i_0_312 (.A1(n_207), .A2(n_0_49__1), .B1(n_0_44__1), .B2(n_206), 
      .ZN(n_0_182));
   AOI221_X1 i_0_313 (.A(n_0_184), .B1(n_205), .B2(n_0_39__1), .C1(n_0_44__1), 
      .C2(n_206), .ZN(n_0_183));
   AOI21_X1 i_0_314 (.A(n_0_185), .B1(n_0_187), .B2(n_0_186), .ZN(n_0_184));
   OAI22_X1 i_0_315 (.A1(n_0_34__1), .A2(n_204), .B1(n_205), .B2(n_0_39__1), 
      .ZN(n_0_185));
   AOI22_X1 i_0_316 (.A1(n_0_34__1), .A2(n_204), .B1(n_203), .B2(n_0_29__1), 
      .ZN(n_0_186));
   OR2_X1 i_0_317 (.A1(n_0_189), .A2(n_0_188), .ZN(n_0_187));
   OAI22_X1 i_0_318 (.A1(n_0_29__1), .A2(n_203), .B1(n_202), .B2(n_0_24__1), 
      .ZN(n_0_188));
   AOI21_X1 i_0_319 (.A(n_0_190), .B1(n_201), .B2(n_0_19__1), .ZN(n_0_189));
   OAI21_X1 i_0_320 (.A(n_0_191), .B1(n_0_193), .B2(n_0_192), .ZN(n_0_190));
   NAND2_X1 i_0_321 (.A1(n_202), .A2(n_0_24__1), .ZN(n_0_191));
   OAI22_X1 i_0_322 (.A1(n_0_19__1), .A2(n_201), .B1(n_200), .B2(n_0_14__1), 
      .ZN(n_0_192));
   AOI221_X1 i_0_323 (.A(n_0_194), .B1(n_199), .B2(n_0_9__1), .C1(n_0_14__1), 
      .C2(n_200), .ZN(n_0_193));
   AOI21_X1 i_0_324 (.A(n_0_195), .B1(n_0_196), .B2(n_109), .ZN(n_0_194));
   OAI22_X1 i_0_325 (.A1(n_0_9__1), .A2(n_199), .B1(n_198), .B2(n_0_4__1), 
      .ZN(n_0_195));
   AOI21_X1 i_0_326 (.A(n_197), .B1(n_198), .B2(n_0_4__1), .ZN(n_0_196));
   NAND2_X1 i_0_327 (.A1(n_77), .A2(n_0_200), .ZN(n_0_197));
   NAND2_X1 i_0_328 (.A1(n_76), .A2(n_0_200), .ZN(n_0_198));
   INV_X1 i_0_329 (.A(n_0_200), .ZN(n_0_199));
   AND2_X1 i_0_330 (.A1(n_65), .A2(n_0_205), .ZN(n_0_200));
   OAI21_X1 i_0_331 (.A(n_0_201), .B1(n_0_277), .B2(n_0), .ZN(n_193));
   NAND2_X1 i_0_332 (.A1(n_0_201), .A2(n_0), .ZN(QuotientVar[15]));
   NAND2_X1 i_0_333 (.A1(n_0_202), .A2(n_0_313), .ZN(n_0_201));
   XNOR2_X1 i_0_334 (.A(n_0_307), .B(Divisor[15]), .ZN(n_0_202));
   AOI21_X1 i_0_335 (.A(Reset), .B1(n_0_262), .B2(n_0_204), .ZN(n_194));
   NOR2_X1 i_0_336 (.A1(Reset), .A2(n_0_203), .ZN(n_195));
   NOR2_X1 i_0_337 (.A1(n_0_286), .A2(Start), .ZN(n_0_203));
   NAND2_X1 i_0_338 (.A1(n_0_205), .A2(n_0_286), .ZN(n_0_204));
   NOR3_X1 i_0_339 (.A1(n_0_206), .A2(n_32), .A3(n_31), .ZN(n_0_205));
   OR3_X1 i_0_340 (.A1(n_0_207), .A2(n_30), .A3(n_29), .ZN(n_0_206));
   INV_X1 i_0_341 (.A(n_0_208), .ZN(n_0_207));
   NOR3_X1 i_0_342 (.A1(n_0_218), .A2(n_0_213), .A3(n_0_209), .ZN(n_0_208));
   NAND3_X1 i_0_343 (.A1(n_0_212), .A2(n_0_211), .A3(n_0_210), .ZN(n_0_209));
   NOR2_X1 i_0_344 (.A1(n_11), .A2(n_12), .ZN(n_0_210));
   NOR2_X1 i_0_345 (.A1(n_9), .A2(n_10), .ZN(n_0_211));
   NOR4_X1 i_0_346 (.A1(n_13), .A2(n_14), .A3(n_15), .A4(n_16), .ZN(n_0_212));
   NAND4_X1 i_0_347 (.A1(n_0_217), .A2(n_0_216), .A3(n_0_215), .A4(n_0_214), 
      .ZN(n_0_213));
   NOR2_X1 i_0_348 (.A1(n_3), .A2(n_4), .ZN(n_0_214));
   NOR2_X1 i_0_349 (.A1(n_1), .A2(n_2), .ZN(n_0_215));
   NOR2_X1 i_0_350 (.A1(n_7), .A2(n_8), .ZN(n_0_216));
   NOR2_X1 i_0_351 (.A1(n_5), .A2(n_6), .ZN(n_0_217));
   NAND3_X1 i_0_352 (.A1(n_0_221), .A2(n_0_220), .A3(n_0_219), .ZN(n_0_218));
   NOR4_X1 i_0_353 (.A1(n_17), .A2(n_18), .A3(n_19), .A4(n_20), .ZN(n_0_219));
   NOR4_X1 i_0_354 (.A1(n_21), .A2(n_22), .A3(n_23), .A4(n_24), .ZN(n_0_220));
   NOR4_X1 i_0_355 (.A1(n_25), .A2(n_26), .A3(n_27), .A4(n_28), .ZN(n_0_221));
   OAI21_X1 i_0_356 (.A(n_0), .B1(n_0_222), .B2(n_0_262), .ZN(n_196));
   AND2_X1 i_0_357 (.A1(n_0_223), .A2(n_0_239), .ZN(n_0_222));
   OAI211_X1 i_0_358 (.A(n_0_245), .B(n_0_224), .C1(n_0_227), .C2(n_0_253), 
      .ZN(n_0_223));
   NOR2_X1 i_0_359 (.A1(n_0_20), .A2(n_0_1), .ZN(n_0_224));
   NOR3_X1 i_0_360 (.A1(n_0_226), .A2(Dividend[12]), .A3(Dividend[13]), .ZN(
      n_0_225));
   OAI21_X1 i_0_361 (.A(n_0_306), .B1(n_0_258), .B2(n_0_255), .ZN(n_0_226));
   NOR3_X1 i_0_362 (.A1(n_0_232), .A2(n_0_228), .A3(n_0_258), .ZN(n_0_227));
   AOI21_X1 i_0_363 (.A(Dividend[14]), .B1(n_0_229), .B2(n_0_256), .ZN(n_0_228));
   OAI211_X1 i_0_364 (.A(n_0_303), .B(n_0_302), .C1(n_0_230), .C2(n_0_255), 
      .ZN(n_0_229));
   AND3_X1 i_0_365 (.A1(n_0_299), .A2(n_0_298), .A3(n_0_231), .ZN(n_0_230));
   OAI211_X1 i_0_366 (.A(n_0_297), .B(n_0_296), .C1(Dividend[3]), .C2(
      Dividend[2]), .ZN(n_0_231));
   NAND2_X1 i_0_367 (.A1(n_0_306), .A2(n_0_233), .ZN(n_0_232));
   OAI21_X1 i_0_368 (.A(n_0_305), .B1(Dividend[12]), .B2(n_0_234), .ZN(n_0_233));
   AOI21_X1 i_0_369 (.A(Dividend[11]), .B1(n_0_302), .B2(n_0_235), .ZN(n_0_234));
   OAI21_X1 i_0_370 (.A(n_0_301), .B1(Dividend[8]), .B2(n_0_236), .ZN(n_0_235));
   AOI21_X1 i_0_371 (.A(Dividend[7]), .B1(n_0_298), .B2(n_0_237), .ZN(n_0_236));
   OAI21_X1 i_0_372 (.A(n_0_297), .B1(Dividend[4]), .B2(n_0_238), .ZN(n_0_237));
   AOI21_X1 i_0_373 (.A(Dividend[3]), .B1(n_0_294), .B2(Dividend[1]), .ZN(
      n_0_238));
   AOI21_X1 i_0_374 (.A(n_0_250), .B1(n_0_245), .B2(n_0_240), .ZN(n_0_239));
   AOI21_X1 i_0_375 (.A(n_0_241), .B1(Divisor[7]), .B2(Divisor[15]), .ZN(n_0_240));
   OR2_X1 i_0_376 (.A1(n_0_242), .A2(Divisor[6]), .ZN(n_0_241));
   OR3_X1 i_0_377 (.A1(n_0_243), .A2(Divisor[4]), .A3(Divisor[5]), .ZN(n_0_242));
   NAND3_X1 i_0_378 (.A1(n_0_244), .A2(n_0_287), .A3(n_0_288), .ZN(n_0_243));
   NOR2_X1 i_0_379 (.A1(Divisor[3]), .A2(Divisor[2]), .ZN(n_0_244));
   NOR3_X1 i_0_380 (.A1(n_0_247), .A2(n_0_246), .A3(Divisor[14]), .ZN(n_0_245));
   OR2_X1 i_0_381 (.A1(Divisor[13]), .A2(Divisor[12]), .ZN(n_0_246));
   NAND2_X1 i_0_382 (.A1(n_0_249), .A2(n_0_248), .ZN(n_0_247));
   NOR2_X1 i_0_383 (.A1(Divisor[9]), .A2(Divisor[8]), .ZN(n_0_248));
   NOR2_X1 i_0_384 (.A1(Divisor[11]), .A2(Divisor[10]), .ZN(n_0_249));
   NOR2_X1 i_0_385 (.A1(n_0_257), .A2(n_0_253), .ZN(n_0_250));
   NAND3_X1 i_0_386 (.A1(n_0_260), .A2(n_0_258), .A3(n_0_254), .ZN(n_0_251));
   NAND4_X1 i_0_387 (.A1(n_0_258), .A2(n_0_300), .A3(n_0_301), .A4(n_0_260), 
      .ZN(n_0_252));
   NAND3_X1 i_0_388 (.A1(n_0_254), .A2(n_0_306), .A3(n_0_256), .ZN(n_0_253));
   INV_X1 i_0_389 (.A(n_0_255), .ZN(n_0_254));
   NAND4_X1 i_0_390 (.A1(n_0_303), .A2(n_0_302), .A3(n_0_301), .A4(n_0_300), 
      .ZN(n_0_255));
   NOR2_X1 i_0_391 (.A1(Dividend[13]), .A2(Dividend[12]), .ZN(n_0_256));
   NAND2_X1 i_0_392 (.A1(n_0_260), .A2(n_0_258), .ZN(n_0_257));
   NOR4_X1 i_0_393 (.A1(Dividend[7]), .A2(Dividend[6]), .A3(Dividend[5]), 
      .A4(Dividend[4]), .ZN(n_0_258));
   NAND3_X1 i_0_394 (.A1(n_0_260), .A2(n_0_296), .A3(n_0_297), .ZN(n_0_259));
   INV_X1 i_0_395 (.A(n_0_261), .ZN(n_0_260));
   NAND4_X1 i_0_396 (.A1(n_0_295), .A2(n_0_294), .A3(n_0_293), .A4(n_0_292), 
      .ZN(n_0_261));
   NAND2_X1 i_0_397 (.A1(Start), .A2(n_0), .ZN(n_0_262));
   AOI21_X1 i_0_398 (.A(n_0_263), .B1(n_126), .B2(n_0_278), .ZN(n_197));
   NOR2_X1 i_0_399 (.A1(n_125), .A2(n_126), .ZN(n_0_263));
   MUX2_X1 i_0_400 (.A(n_124), .B(addOut[1]), .S(n_126), .Z(n_198));
   MUX2_X1 i_0_401 (.A(n_123), .B(addOut[2]), .S(n_126), .Z(n_199));
   MUX2_X1 i_0_402 (.A(n_122), .B(addOut[3]), .S(n_126), .Z(n_200));
   AOI21_X1 i_0_403 (.A(n_0_264), .B1(n_126), .B2(n_0_279), .ZN(n_201));
   NOR2_X1 i_0_404 (.A1(n_121), .A2(n_126), .ZN(n_0_264));
   AOI21_X1 i_0_405 (.A(n_0_265), .B1(n_126), .B2(n_0_280), .ZN(n_202));
   NOR2_X1 i_0_406 (.A1(n_120), .A2(n_126), .ZN(n_0_265));
   MUX2_X1 i_0_407 (.A(n_119), .B(addOut[6]), .S(n_126), .Z(n_203));
   MUX2_X1 i_0_408 (.A(n_118), .B(addOut[7]), .S(n_126), .Z(n_204));
   AOI21_X1 i_0_409 (.A(n_0_266), .B1(n_126), .B2(n_0_281), .ZN(n_205));
   NOR2_X1 i_0_410 (.A1(n_117), .A2(n_126), .ZN(n_0_266));
   AOI21_X1 i_0_411 (.A(n_0_267), .B1(n_126), .B2(n_0_282), .ZN(n_206));
   NOR2_X1 i_0_412 (.A1(n_116), .A2(n_126), .ZN(n_0_267));
   MUX2_X1 i_0_413 (.A(n_115), .B(addOut[10]), .S(n_126), .Z(n_207));
   MUX2_X1 i_0_414 (.A(n_114), .B(addOut[11]), .S(n_126), .Z(n_208));
   AOI21_X1 i_0_415 (.A(n_0_268), .B1(n_126), .B2(n_0_283), .ZN(n_209));
   NOR2_X1 i_0_416 (.A1(n_113), .A2(n_126), .ZN(n_0_268));
   MUX2_X1 i_0_417 (.A(n_112), .B(addOut[13]), .S(n_126), .Z(n_210));
   MUX2_X1 i_0_418 (.A(n_111), .B(addOut[14]), .S(n_126), .Z(n_211));
   INV_X1 i_0_419 (.A(n_0_269), .ZN(n_212));
   OAI21_X1 i_0_420 (.A(n_0_270), .B1(n_126), .B2(n_110), .ZN(n_0_269));
   NAND2_X1 i_0_421 (.A1(n_0_284), .A2(n_126), .ZN(n_0_270));
   INV_X1 i_0_422 (.A(n_35), .ZN(n_0_271));
   INV_X1 i_0_423 (.A(n_37), .ZN(n_0_272));
   INV_X1 i_0_424 (.A(n_79), .ZN(n_0_273));
   INV_X1 i_0_425 (.A(n_74), .ZN(n_0_274));
   INV_X1 i_0_426 (.A(n_71), .ZN(n_0_275));
   INV_X1 i_0_427 (.A(n_68), .ZN(n_0_276));
   INV_X1 i_0_428 (.A(n_65), .ZN(n_0_277));
   INV_X1 i_0_429 (.A(addOut[0]), .ZN(n_0_278));
   INV_X1 i_0_430 (.A(addOut[4]), .ZN(n_0_279));
   INV_X1 i_0_431 (.A(addOut[5]), .ZN(n_0_280));
   INV_X1 i_0_432 (.A(addOut[8]), .ZN(n_0_281));
   INV_X1 i_0_433 (.A(addOut[9]), .ZN(n_0_282));
   INV_X1 i_0_434 (.A(addOut[12]), .ZN(n_0_283));
   INV_X1 i_0_435 (.A(addOut[15]), .ZN(n_0_284));
   INV_X1 i_0_436 (.A(Reset), .ZN(n_0_285));
   INV_X1 i_0_437 (.A(n_0), .ZN(n_0_286));
   INV_X1 i_0_438 (.A(Divisor[0]), .ZN(n_0_287));
   INV_X1 i_0_439 (.A(Divisor[1]), .ZN(n_0_288));
   INV_X1 i_0_440 (.A(Divisor[2]), .ZN(n_0_289));
   INV_X1 i_0_441 (.A(Divisor[10]), .ZN(n_0_290));
   INV_X1 i_0_442 (.A(Divisor[15]), .ZN(n_0_291));
   INV_X1 i_0_443 (.A(Dividend[0]), .ZN(n_0_292));
   INV_X1 i_0_444 (.A(Dividend[1]), .ZN(n_0_293));
   INV_X1 i_0_445 (.A(Dividend[2]), .ZN(n_0_294));
   INV_X1 i_0_446 (.A(Dividend[3]), .ZN(n_0_295));
   INV_X1 i_0_447 (.A(Dividend[4]), .ZN(n_0_296));
   INV_X1 i_0_448 (.A(Dividend[5]), .ZN(n_0_297));
   INV_X1 i_0_449 (.A(Dividend[6]), .ZN(n_0_298));
   INV_X1 i_0_450 (.A(Dividend[7]), .ZN(n_0_299));
   INV_X1 i_0_451 (.A(Dividend[8]), .ZN(n_0_300));
   INV_X1 i_0_452 (.A(Dividend[9]), .ZN(n_0_301));
   INV_X1 i_0_453 (.A(Dividend[10]), .ZN(n_0_302));
   INV_X1 i_0_454 (.A(Dividend[11]), .ZN(n_0_303));
   INV_X1 i_0_455 (.A(Dividend[12]), .ZN(n_0_304));
   INV_X1 i_0_456 (.A(Dividend[13]), .ZN(n_0_305));
   INV_X1 i_0_457 (.A(Dividend[14]), .ZN(n_0_306));
   INV_X1 i_0_458 (.A(Dividend[15]), .ZN(n_0_307));
   INV_X1 i_0_459 (.A(n_30), .ZN(n_0_308));
   INV_X1 i_0_460 (.A(n_109), .ZN(n_213));
   INV_X1 i_0_461 (.A(n_108), .ZN(n_0_4__1));
   INV_X1 i_0_462 (.A(n_107), .ZN(n_0_9__1));
   INV_X1 i_0_463 (.A(n_106), .ZN(n_0_14__1));
   INV_X1 i_0_464 (.A(n_105), .ZN(n_0_19__1));
   INV_X1 i_0_465 (.A(n_104), .ZN(n_0_24__1));
   INV_X1 i_0_466 (.A(n_103), .ZN(n_0_29__1));
   INV_X1 i_0_467 (.A(n_102), .ZN(n_0_34__1));
   INV_X1 i_0_468 (.A(n_101), .ZN(n_0_39__1));
   INV_X1 i_0_469 (.A(n_100), .ZN(n_0_44__1));
   INV_X1 i_0_470 (.A(n_99), .ZN(n_0_49__1));
   INV_X1 i_0_471 (.A(n_98), .ZN(n_0_54__1));
   INV_X1 i_0_472 (.A(n_97), .ZN(n_0_59__1));
   INV_X1 i_0_473 (.A(n_96), .ZN(n_0_64__1));
   INV_X1 i_0_474 (.A(n_95), .ZN(n_0_69__1));
   INV_X1 i_0_475 (.A(n_94), .ZN(n_0_74__1));
   INV_X1 i_0_476 (.A(n_92), .ZN(n_0_309));
   INV_X1 i_0_477 (.A(n_91), .ZN(n_0_310));
   INV_X1 i_0_478 (.A(n_89), .ZN(n_0_311));
   INV_X1 i_0_479 (.A(n_88), .ZN(n_0_312));
   INV_X1 i_0_480 (.A(n_0_262), .ZN(n_0_313));
endmodule

module StepAlgo(h_in, L, e, test, reset, CLK, EN, Done, h_new);
   input [15:0]h_in;
   input [15:0]L;
   input [15:0]e;
   input [15:0]test;
   input reset;
   input CLK;
   input EN;
   output Done;
   output [15:0]h_new;

   wire Q2;
   wire Q1;
   wire DoneSignal;
   wire [15:0]Division_output;
   wire L1;
   wire n_0_0;

   flipflop__2_64 F2 (.D(EN), .load(Q1), .Clk(CLK), .Q(Q2), .rst());
   flipflop F (.D(EN), .load(L1), .Clk(CLK), .Q(Q1), .rst(Q2));
   fixed_division D1 (.Dividend(test), .Divisor(e), .Reset(reset), .clk(), 
      .Start(Q1), .Quotient(Division_output), .ERR(), .Done(DoneSignal), 
      .OverFlow());
   TBUF_X1 i_0_1 (.A(Division_output[0]), .EN(n_0_0), .Z(h_new[0]));
   TBUF_X1 i_0_2 (.A(Division_output[1]), .EN(n_0_0), .Z(h_new[1]));
   TBUF_X1 i_0_3 (.A(Division_output[2]), .EN(n_0_0), .Z(h_new[2]));
   TBUF_X1 i_0_4 (.A(Division_output[3]), .EN(n_0_0), .Z(h_new[3]));
   TBUF_X1 i_0_5 (.A(Division_output[4]), .EN(n_0_0), .Z(h_new[4]));
   TBUF_X1 i_0_6 (.A(Division_output[5]), .EN(n_0_0), .Z(h_new[5]));
   TBUF_X1 i_0_7 (.A(Division_output[6]), .EN(n_0_0), .Z(h_new[6]));
   TBUF_X1 i_0_8 (.A(Division_output[7]), .EN(n_0_0), .Z(h_new[7]));
   TBUF_X1 i_0_9 (.A(Division_output[8]), .EN(n_0_0), .Z(h_new[8]));
   TBUF_X1 i_0_10 (.A(Division_output[9]), .EN(n_0_0), .Z(h_new[9]));
   TBUF_X1 i_0_11 (.A(Division_output[10]), .EN(n_0_0), .Z(h_new[10]));
   TBUF_X1 i_0_12 (.A(Division_output[11]), .EN(n_0_0), .Z(h_new[11]));
   TBUF_X1 i_0_13 (.A(Division_output[12]), .EN(n_0_0), .Z(h_new[12]));
   TBUF_X1 i_0_14 (.A(Division_output[13]), .EN(n_0_0), .Z(h_new[13]));
   TBUF_X1 i_0_15 (.A(Division_output[14]), .EN(n_0_0), .Z(h_new[14]));
   TBUF_X1 i_0_16 (.A(Division_output[15]), .EN(n_0_0), .Z(h_new[15]));
   INV_X1 i_0_0_0 (.A(reset), .ZN(L1));
   AND2_X1 i_0_17_0 (.A1(DoneSignal), .A2(EN), .ZN(Done));
   NOR2_X1 i_0_17_1 (.A1(DoneSignal), .A2(EN), .ZN(n_0_0));
endmodule
