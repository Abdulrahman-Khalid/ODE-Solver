/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 23:33:54 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 508608438 */

module Partial_Full_Adder__0_66(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   INV_X1 i_3 (.A(P), .ZN(S));
   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_70(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_74(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_78(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_82(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_86(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_90(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_94(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_98(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_102(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_106(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_110(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_114(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_118(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_122(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire G;
   wire P;
   wire c15;
   wire n_0_0;
   wire c14;
   wire n_0_1;
   wire c13;
   wire n_0_2;
   wire c12;
   wire n_0_3;
   wire c11;
   wire n_0_4;
   wire c10;
   wire n_0_5;
   wire c9;
   wire n_0_6;
   wire c8;
   wire n_0_7;
   wire c7;
   wire n_0_8;
   wire c6;
   wire n_0_9;
   wire c5;
   wire n_0_10;
   wire c4;
   wire n_0_11;
   wire c3;
   wire n_0_12;
   wire c2;
   wire n_0_13;
   wire c1;

   Partial_Full_Adder__0_66 PFA1 (.A(A[0]), .B(B[0]), .Cin(), .S(S[0]), .P(P), 
      .G(G));
   Partial_Full_Adder__0_70 PFA2 (.A(A[1]), .B(B[1]), .Cin(c1), .S(S[1]), 
      .P(n_1), .G(n_0));
   Partial_Full_Adder__0_74 PFA3 (.A(A[2]), .B(B[2]), .Cin(c2), .S(S[2]), 
      .P(n_3), .G(n_2));
   Partial_Full_Adder__0_78 PFA4 (.A(A[3]), .B(B[3]), .Cin(c3), .S(S[3]), 
      .P(n_5), .G(n_4));
   Partial_Full_Adder__0_82 PFA5 (.A(A[4]), .B(B[4]), .Cin(c4), .S(S[4]), 
      .P(n_7), .G(n_6));
   Partial_Full_Adder__0_86 PFA6 (.A(A[5]), .B(B[5]), .Cin(c5), .S(S[5]), 
      .P(n_9), .G(n_8));
   Partial_Full_Adder__0_90 PFA7 (.A(A[6]), .B(B[6]), .Cin(c6), .S(S[6]), 
      .P(n_11), .G(n_10));
   Partial_Full_Adder__0_94 PFA8 (.A(A[7]), .B(B[7]), .Cin(c7), .S(S[7]), 
      .P(n_13), .G(n_12));
   Partial_Full_Adder__0_98 PFA9 (.A(A[8]), .B(B[8]), .Cin(c8), .S(S[8]), 
      .P(n_15), .G(n_14));
   Partial_Full_Adder__0_102 PFA10 (.A(A[9]), .B(B[9]), .Cin(c9), .S(S[9]), 
      .P(n_17), .G(n_16));
   Partial_Full_Adder__0_106 PFA11 (.A(A[10]), .B(B[10]), .Cin(c10), .S(S[10]), 
      .P(n_19), .G(n_18));
   Partial_Full_Adder__0_110 PFA12 (.A(A[11]), .B(B[11]), .Cin(c11), .S(S[11]), 
      .P(n_21), .G(n_20));
   Partial_Full_Adder__0_114 PFA13 (.A(A[12]), .B(B[12]), .Cin(c12), .S(S[12]), 
      .P(n_23), .G(n_22));
   Partial_Full_Adder__0_118 PFA14 (.A(A[13]), .B(B[13]), .Cin(c13), .S(S[13]), 
      .P(n_25), .G(n_24));
   Partial_Full_Adder__0_122 PFA15 (.A(A[14]), .B(B[14]), .Cin(c14), .S(S[14]), 
      .P(n_27), .G(n_26));
   Partial_Full_Adder PFA16 (.A(A[15]), .B(B[15]), .Cin(c15), .S(S[15]), .P(), 
      .G());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(c15));
   AOI21_X1 i_0_1 (.A(n_26), .B1(n_27), .B2(c14), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(c14));
   AOI21_X1 i_0_3 (.A(n_24), .B1(n_25), .B2(c13), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(c13));
   AOI21_X1 i_0_5 (.A(n_22), .B1(n_23), .B2(c12), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(c12));
   AOI21_X1 i_0_7 (.A(n_20), .B1(n_21), .B2(c11), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(c11));
   AOI21_X1 i_0_9 (.A(n_18), .B1(n_19), .B2(c10), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(c10));
   AOI21_X1 i_0_11 (.A(n_16), .B1(n_17), .B2(c9), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(c9));
   AOI21_X1 i_0_13 (.A(n_14), .B1(n_15), .B2(c8), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(c8));
   AOI21_X1 i_0_15 (.A(n_12), .B1(n_13), .B2(c7), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(c7));
   AOI21_X1 i_0_17 (.A(n_10), .B1(n_11), .B2(c6), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(c6));
   AOI21_X1 i_0_19 (.A(n_8), .B1(n_9), .B2(c5), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(c5));
   AOI21_X1 i_0_21 (.A(n_6), .B1(n_7), .B2(c4), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(c4));
   AOI21_X1 i_0_23 (.A(n_4), .B1(n_5), .B2(c3), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(c3));
   AOI21_X1 i_0_25 (.A(n_2), .B1(n_3), .B2(c2), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(c2));
   AOI21_X1 i_0_27 (.A(n_0), .B1(n_1), .B2(c1), .ZN(n_0_13));
   OR2_X1 i_0_28 (.A1(P), .A2(G), .ZN(c1));
endmodule

module datapath__0_49(Index, p_0);
   input [31:0]Index;
   output [31:0]p_0;

   XNOR2_X1 i_1 (.A(Index[1]), .B(Index[0]), .ZN(p_0[1]));
   OR2_X1 i_2 (.A1(Index[1]), .A2(Index[0]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(Index[2]), .B(n_0), .ZN(p_0[2]));
   OR2_X1 i_4 (.A1(Index[2]), .A2(n_0), .ZN(n_1));
   XNOR2_X1 i_5 (.A(Index[3]), .B(n_1), .ZN(p_0[3]));
   OR2_X1 i_6 (.A1(Index[3]), .A2(n_1), .ZN(n_2));
   XNOR2_X1 i_7 (.A(Index[4]), .B(n_2), .ZN(p_0[4]));
   OR2_X1 i_8 (.A1(Index[4]), .A2(n_2), .ZN(n_3));
   XNOR2_X1 i_9 (.A(Index[5]), .B(n_3), .ZN(p_0[5]));
   OR2_X1 i_10 (.A1(Index[5]), .A2(n_3), .ZN(n_4));
   XNOR2_X1 i_11 (.A(Index[6]), .B(n_4), .ZN(p_0[6]));
   OR2_X1 i_12 (.A1(Index[6]), .A2(n_4), .ZN(n_5));
   XNOR2_X1 i_13 (.A(Index[7]), .B(n_5), .ZN(p_0[7]));
   OR2_X1 i_14 (.A1(Index[7]), .A2(n_5), .ZN(n_6));
   XNOR2_X1 i_15 (.A(Index[8]), .B(n_6), .ZN(p_0[8]));
   OR2_X1 i_16 (.A1(Index[8]), .A2(n_6), .ZN(n_7));
   XNOR2_X1 i_17 (.A(Index[9]), .B(n_7), .ZN(p_0[9]));
   OR2_X1 i_18 (.A1(Index[9]), .A2(n_7), .ZN(n_8));
   XNOR2_X1 i_19 (.A(Index[10]), .B(n_8), .ZN(p_0[10]));
   OR2_X1 i_20 (.A1(Index[10]), .A2(n_8), .ZN(n_9));
   XNOR2_X1 i_21 (.A(Index[11]), .B(n_9), .ZN(p_0[11]));
   OR2_X1 i_22 (.A1(Index[11]), .A2(n_9), .ZN(n_10));
   XNOR2_X1 i_23 (.A(Index[12]), .B(n_10), .ZN(p_0[12]));
   OR2_X1 i_24 (.A1(Index[12]), .A2(n_10), .ZN(n_11));
   XNOR2_X1 i_25 (.A(Index[13]), .B(n_11), .ZN(p_0[13]));
   OR2_X1 i_26 (.A1(Index[13]), .A2(n_11), .ZN(n_12));
   XNOR2_X1 i_27 (.A(Index[14]), .B(n_12), .ZN(p_0[14]));
   OR2_X1 i_28 (.A1(Index[14]), .A2(n_12), .ZN(n_13));
   XNOR2_X1 i_29 (.A(Index[15]), .B(n_13), .ZN(p_0[15]));
   OR2_X1 i_30 (.A1(Index[15]), .A2(n_13), .ZN(n_14));
   XNOR2_X1 i_31 (.A(Index[16]), .B(n_14), .ZN(p_0[16]));
   OR2_X1 i_32 (.A1(Index[16]), .A2(n_14), .ZN(n_15));
   XNOR2_X1 i_33 (.A(Index[17]), .B(n_15), .ZN(p_0[17]));
   OR2_X1 i_34 (.A1(Index[17]), .A2(n_15), .ZN(n_16));
   XNOR2_X1 i_35 (.A(Index[18]), .B(n_16), .ZN(p_0[18]));
   OR2_X1 i_36 (.A1(Index[18]), .A2(n_16), .ZN(n_17));
   XNOR2_X1 i_37 (.A(Index[19]), .B(n_17), .ZN(p_0[19]));
   OR2_X1 i_38 (.A1(Index[19]), .A2(n_17), .ZN(n_18));
   XNOR2_X1 i_39 (.A(Index[20]), .B(n_18), .ZN(p_0[20]));
   OR2_X1 i_40 (.A1(Index[20]), .A2(n_18), .ZN(n_19));
   XNOR2_X1 i_41 (.A(Index[21]), .B(n_19), .ZN(p_0[21]));
   OR2_X1 i_42 (.A1(Index[21]), .A2(n_19), .ZN(n_20));
   XNOR2_X1 i_43 (.A(Index[22]), .B(n_20), .ZN(p_0[22]));
   OR2_X1 i_44 (.A1(Index[22]), .A2(n_20), .ZN(n_21));
   XNOR2_X1 i_45 (.A(Index[23]), .B(n_21), .ZN(p_0[23]));
   OR2_X1 i_46 (.A1(Index[23]), .A2(n_21), .ZN(n_22));
   XNOR2_X1 i_47 (.A(Index[24]), .B(n_22), .ZN(p_0[24]));
   OR2_X1 i_48 (.A1(Index[24]), .A2(n_22), .ZN(n_23));
   XNOR2_X1 i_49 (.A(Index[25]), .B(n_23), .ZN(p_0[25]));
   OR2_X1 i_50 (.A1(Index[25]), .A2(n_23), .ZN(n_24));
   XNOR2_X1 i_51 (.A(Index[26]), .B(n_24), .ZN(p_0[26]));
   OR2_X1 i_52 (.A1(Index[26]), .A2(n_24), .ZN(n_25));
   XNOR2_X1 i_53 (.A(Index[27]), .B(n_25), .ZN(p_0[27]));
   OR2_X1 i_54 (.A1(Index[27]), .A2(n_25), .ZN(n_26));
   XNOR2_X1 i_55 (.A(Index[28]), .B(n_26), .ZN(p_0[28]));
   OR2_X1 i_56 (.A1(Index[28]), .A2(n_26), .ZN(n_27));
   XNOR2_X1 i_57 (.A(Index[29]), .B(n_27), .ZN(p_0[29]));
   OR2_X1 i_58 (.A1(Index[29]), .A2(n_27), .ZN(n_28));
   XNOR2_X1 i_59 (.A(Index[30]), .B(n_28), .ZN(p_0[30]));
   OR2_X1 i_60 (.A1(Index[30]), .A2(n_28), .ZN(n_29));
   XNOR2_X1 i_61 (.A(Index[31]), .B(n_29), .ZN(p_0[31]));
endmodule

module fixed_division(Dividend, Divisor, rst, clk, Start, Quotient, ERR, Done, 
      OverFlow);
   input [15:0]Dividend;
   input [15:0]Divisor;
   input rst;
   input clk;
   input Start;
   output [15:0]Quotient;
   output ERR;
   output Done;
   output OverFlow;

   wire [15:0]addOut;
   wire n_0_1;
   wire n_0_25;
   wire [15:0]add2;
   wire [15:0]add1;
   wire n_0_2;
   wire [31:0]Index;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire [15:0]QuotientVar;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire [15:0]Dividend2;
   wire n_0_0;
   wire n_0_64;
   wire FIRST_ONE;
   wire n_0_65;
   wire n_0_159;
   wire n_0_142;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_16;
   wire n_0_0_2;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_3;
   wire n_0_0_13;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_66;
   wire n_0_0_27;
   wire n_0_69;
   wire n_0_68;
   wire n_0_70;
   wire n_0_71;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_72;
   wire n_0_0_30;
   wire n_0_73;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_74;
   wire n_0_0_34;
   wire n_0_75;
   wire n_0_0_35;
   wire n_0_76;
   wire n_0_0_36;
   wire n_0_77;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_78;
   wire n_0_0_44;
   wire n_0_79;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_80;
   wire n_0_0_47;
   wire n_0_81;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_82;
   wire n_0_0_52;
   wire n_0_83;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_84;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_0_59;
   wire n_0_101;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_102;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_103;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_104;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_105;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_106;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_107;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_108;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_109;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_110;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_111;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_112;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_113;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_114;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_0_106;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_130;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_0_107;
   wire n_0_67;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_0_108;
   wire n_0_201;
   wire n_0_0_109;
   wire n_0_202;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_203;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_204;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_205;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_206;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_207;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_208;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_209;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_210;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_211;
   wire n_0_0_128;
   wire n_0_212;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_213;
   wire n_0_0_131;
   wire n_0_214;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_215;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_216;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_217;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_218;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_219;
   wire n_0_0_272;
   wire n_0_220;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_222;
   wire n_0_221;

   Carry_Look_Ahead u1 (.A(add1), .B(add2), .Cin(), .S(addOut));
   DFF_X1 Done_reg (.D(n_0_1), .CK(clk), .Q(Done), .QN());
   MUX2_X1 Done_reg_enable_mux_0 (.A(Done), .B(n_0_218), .S(n_0_217), .Z(n_0_1));
   CLKGATETST_X1 clk_gate_Quotient_reg (.CK(clk), .E(n_0_199), .SE(1'b0), 
      .GCK(n_0_25));
   DFF_X1 \Quotient_reg[15]  (.D(n_0_215), .CK(n_0_25), .Q(Quotient[15]), .QN());
   DFF_X1 \Quotient_reg[14]  (.D(n_0_214), .CK(n_0_25), .Q(Quotient[14]), .QN());
   DFF_X1 \Quotient_reg[13]  (.D(n_0_213), .CK(n_0_25), .Q(Quotient[13]), .QN());
   DFF_X1 \Quotient_reg[12]  (.D(n_0_212), .CK(n_0_25), .Q(Quotient[12]), .QN());
   DFF_X1 \Quotient_reg[11]  (.D(n_0_211), .CK(n_0_25), .Q(Quotient[11]), .QN());
   DFF_X1 \Quotient_reg[10]  (.D(n_0_210), .CK(n_0_25), .Q(Quotient[10]), .QN());
   DFF_X1 \Quotient_reg[9]  (.D(n_0_209), .CK(n_0_25), .Q(Quotient[9]), .QN());
   DFF_X1 \Quotient_reg[8]  (.D(n_0_208), .CK(n_0_25), .Q(Quotient[8]), .QN());
   DFF_X1 \Quotient_reg[7]  (.D(n_0_207), .CK(n_0_25), .Q(Quotient[7]), .QN());
   DFF_X1 \Quotient_reg[6]  (.D(n_0_206), .CK(n_0_25), .Q(Quotient[6]), .QN());
   DFF_X1 \Quotient_reg[5]  (.D(n_0_205), .CK(n_0_25), .Q(Quotient[5]), .QN());
   DFF_X1 \Quotient_reg[4]  (.D(n_0_204), .CK(n_0_25), .Q(Quotient[4]), .QN());
   DFF_X1 \Quotient_reg[3]  (.D(n_0_203), .CK(n_0_25), .Q(Quotient[3]), .QN());
   DFF_X1 \Quotient_reg[2]  (.D(n_0_202), .CK(n_0_25), .Q(Quotient[2]), .QN());
   DFF_X1 \Quotient_reg[1]  (.D(n_0_201), .CK(n_0_25), .Q(Quotient[1]), .QN());
   DFF_X1 \Quotient_reg[0]  (.D(n_0_200), .CK(n_0_25), .Q(Quotient[0]), .QN());
   DFF_X1 \add2_reg[15]  (.D(n_0_198), .CK(n_0_142), .Q(add2[15]), .QN());
   DFF_X1 \add2_reg[14]  (.D(n_0_197), .CK(n_0_142), .Q(add2[14]), .QN());
   DFF_X1 \add2_reg[13]  (.D(n_0_196), .CK(n_0_142), .Q(add2[13]), .QN());
   DFF_X1 \add2_reg[12]  (.D(n_0_195), .CK(n_0_142), .Q(add2[12]), .QN());
   DFF_X1 \add2_reg[11]  (.D(n_0_194), .CK(n_0_142), .Q(add2[11]), .QN());
   DFF_X1 \add2_reg[10]  (.D(n_0_193), .CK(n_0_142), .Q(add2[10]), .QN());
   DFF_X1 \add2_reg[9]  (.D(n_0_192), .CK(n_0_142), .Q(add2[9]), .QN());
   DFF_X1 \add2_reg[8]  (.D(n_0_191), .CK(n_0_142), .Q(add2[8]), .QN());
   DFF_X1 \add2_reg[7]  (.D(n_0_190), .CK(n_0_142), .Q(add2[7]), .QN());
   DFF_X1 \add2_reg[6]  (.D(n_0_189), .CK(n_0_142), .Q(add2[6]), .QN());
   DFF_X1 \add2_reg[5]  (.D(n_0_188), .CK(n_0_142), .Q(add2[5]), .QN());
   DFF_X1 \add2_reg[4]  (.D(n_0_187), .CK(n_0_142), .Q(add2[4]), .QN());
   DFF_X1 \add2_reg[3]  (.D(n_0_186), .CK(n_0_142), .Q(add2[3]), .QN());
   DFF_X1 \add2_reg[2]  (.D(n_0_185), .CK(n_0_142), .Q(add2[2]), .QN());
   DFF_X1 \add2_reg[1]  (.D(n_0_184), .CK(n_0_142), .Q(add2[1]), .QN());
   DFF_X1 \add2_reg[0]  (.D(n_0_183), .CK(n_0_142), .Q(add2[0]), .QN());
   DFF_X1 \add1_reg[15]  (.D(n_0_181), .CK(n_0_142), .Q(add1[15]), .QN());
   DFF_X1 \add1_reg[14]  (.D(n_0_180), .CK(n_0_142), .Q(add1[14]), .QN());
   DFF_X1 \add1_reg[13]  (.D(n_0_179), .CK(n_0_142), .Q(add1[13]), .QN());
   DFF_X1 \add1_reg[12]  (.D(n_0_178), .CK(n_0_142), .Q(add1[12]), .QN());
   DFF_X1 \add1_reg[11]  (.D(n_0_177), .CK(n_0_142), .Q(add1[11]), .QN());
   DFF_X1 \add1_reg[10]  (.D(n_0_176), .CK(n_0_142), .Q(add1[10]), .QN());
   DFF_X1 \add1_reg[9]  (.D(n_0_175), .CK(n_0_142), .Q(add1[9]), .QN());
   DFF_X1 \add1_reg[8]  (.D(n_0_174), .CK(n_0_142), .Q(add1[8]), .QN());
   DFF_X1 \add1_reg[7]  (.D(n_0_173), .CK(n_0_142), .Q(add1[7]), .QN());
   DFF_X1 \add1_reg[6]  (.D(n_0_172), .CK(n_0_142), .Q(add1[6]), .QN());
   DFF_X1 \add1_reg[5]  (.D(n_0_171), .CK(n_0_142), .Q(add1[5]), .QN());
   DFF_X1 \add1_reg[4]  (.D(n_0_170), .CK(n_0_142), .Q(add1[4]), .QN());
   DFF_X1 \add1_reg[3]  (.D(n_0_169), .CK(n_0_142), .Q(add1[3]), .QN());
   DFF_X1 \add1_reg[2]  (.D(n_0_168), .CK(n_0_142), .Q(add1[2]), .QN());
   DFF_X1 \add1_reg[1]  (.D(n_0_167), .CK(n_0_142), .Q(add1[1]), .QN());
   DFF_X1 \add1_reg[0]  (.D(n_0_166), .CK(n_0_142), .Q(add1[0]), .QN());
   DFF_X1 Done_bit_reg (.D(n_0_165), .CK(n_0_159), .Q(n_0_2), .QN());
   DFF_X1 \Index_reg[31]  (.D(n_0_164), .CK(n_0_159), .Q(Index[31]), .QN());
   DFF_X1 \Index_reg[30]  (.D(n_0_163), .CK(n_0_159), .Q(Index[30]), .QN());
   DFF_X1 \Index_reg[29]  (.D(n_0_162), .CK(n_0_159), .Q(Index[29]), .QN());
   DFF_X1 \Index_reg[28]  (.D(n_0_161), .CK(n_0_159), .Q(Index[28]), .QN());
   DFF_X1 \Index_reg[27]  (.D(n_0_160), .CK(n_0_159), .Q(Index[27]), .QN());
   DFF_X1 \Index_reg[26]  (.D(n_0_158), .CK(n_0_159), .Q(Index[26]), .QN());
   DFF_X1 \Index_reg[25]  (.D(n_0_157), .CK(n_0_159), .Q(Index[25]), .QN());
   DFF_X1 \Index_reg[24]  (.D(n_0_156), .CK(n_0_159), .Q(Index[24]), .QN());
   DFF_X1 \Index_reg[23]  (.D(n_0_155), .CK(n_0_159), .Q(Index[23]), .QN());
   DFF_X1 \Index_reg[22]  (.D(n_0_154), .CK(n_0_159), .Q(Index[22]), .QN());
   DFF_X1 \Index_reg[21]  (.D(n_0_153), .CK(n_0_159), .Q(Index[21]), .QN());
   DFF_X1 \Index_reg[20]  (.D(n_0_152), .CK(n_0_159), .Q(Index[20]), .QN());
   DFF_X1 \Index_reg[19]  (.D(n_0_151), .CK(n_0_159), .Q(Index[19]), .QN());
   DFF_X1 \Index_reg[18]  (.D(n_0_150), .CK(n_0_159), .Q(Index[18]), .QN());
   DFF_X1 \Index_reg[17]  (.D(n_0_149), .CK(n_0_159), .Q(Index[17]), .QN());
   DFF_X1 \Index_reg[16]  (.D(n_0_148), .CK(n_0_159), .Q(Index[16]), .QN());
   DFF_X1 \Index_reg[15]  (.D(n_0_147), .CK(n_0_159), .Q(Index[15]), .QN());
   DFF_X1 \Index_reg[14]  (.D(n_0_146), .CK(n_0_159), .Q(Index[14]), .QN());
   DFF_X1 \Index_reg[13]  (.D(n_0_145), .CK(n_0_159), .Q(Index[13]), .QN());
   DFF_X1 \Index_reg[12]  (.D(n_0_144), .CK(n_0_159), .Q(Index[12]), .QN());
   DFF_X1 \Index_reg[11]  (.D(n_0_143), .CK(n_0_159), .Q(Index[11]), .QN());
   DFF_X1 \Index_reg[10]  (.D(n_0_141), .CK(n_0_159), .Q(Index[10]), .QN());
   DFF_X1 \Index_reg[9]  (.D(n_0_140), .CK(n_0_159), .Q(Index[9]), .QN());
   DFF_X1 \Index_reg[8]  (.D(n_0_139), .CK(n_0_159), .Q(Index[8]), .QN());
   DFF_X1 \Index_reg[7]  (.D(n_0_138), .CK(n_0_159), .Q(Index[7]), .QN());
   DFF_X1 \Index_reg[6]  (.D(n_0_137), .CK(n_0_159), .Q(Index[6]), .QN());
   DFF_X1 \Index_reg[5]  (.D(n_0_136), .CK(n_0_159), .Q(Index[5]), .QN());
   DFF_X1 \Index_reg[4]  (.D(n_0_135), .CK(n_0_159), .Q(Index[4]), .QN());
   DFF_X1 \Index_reg[3]  (.D(n_0_134), .CK(n_0_159), .Q(Index[3]), .QN());
   DFF_X1 \Index_reg[2]  (.D(n_0_133), .CK(n_0_159), .Q(Index[2]), .QN());
   DFF_X1 \Index_reg[1]  (.D(n_0_132), .CK(n_0_159), .Q(Index[1]), .QN());
   DFF_X1 \Index_reg[0]  (.D(n_0_131), .CK(n_0_159), .Q(Index[0]), .QN());
   datapath__0_49 i_0_32 (.Index(Index), .p_0({n_0_34, n_0_33, n_0_32, n_0_31, 
      n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_24, n_0_23, n_0_22, n_0_21, 
      n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, uc_0}));
   DFF_X1 \QuotientVar_reg[15]  (.D(n_0_215), .CK(n_0_159), .Q(QuotientVar[15]), 
      .QN());
   DFF_X1 \QuotientVar_reg[14]  (.D(n_0_129), .CK(n_0_159), .Q(QuotientVar[14]), 
      .QN());
   DFF_X1 \QuotientVar_reg[13]  (.D(n_0_128), .CK(n_0_159), .Q(QuotientVar[13]), 
      .QN());
   DFF_X1 \QuotientVar_reg[12]  (.D(n_0_127), .CK(n_0_159), .Q(QuotientVar[12]), 
      .QN());
   DFF_X1 \QuotientVar_reg[11]  (.D(n_0_126), .CK(n_0_159), .Q(QuotientVar[11]), 
      .QN());
   DFF_X1 \QuotientVar_reg[10]  (.D(n_0_125), .CK(n_0_159), .Q(QuotientVar[10]), 
      .QN());
   DFF_X1 \QuotientVar_reg[9]  (.D(n_0_124), .CK(n_0_159), .Q(QuotientVar[9]), 
      .QN());
   DFF_X1 \QuotientVar_reg[8]  (.D(n_0_123), .CK(n_0_159), .Q(QuotientVar[8]), 
      .QN());
   DFF_X1 \QuotientVar_reg[7]  (.D(n_0_122), .CK(n_0_159), .Q(QuotientVar[7]), 
      .QN());
   DFF_X1 \QuotientVar_reg[6]  (.D(n_0_121), .CK(n_0_159), .Q(QuotientVar[6]), 
      .QN());
   DFF_X1 \QuotientVar_reg[5]  (.D(n_0_120), .CK(n_0_159), .Q(QuotientVar[5]), 
      .QN());
   DFF_X1 \QuotientVar_reg[4]  (.D(n_0_119), .CK(n_0_159), .Q(QuotientVar[4]), 
      .QN());
   DFF_X1 \QuotientVar_reg[3]  (.D(n_0_118), .CK(n_0_159), .Q(QuotientVar[3]), 
      .QN());
   DFF_X1 \QuotientVar_reg[2]  (.D(n_0_117), .CK(n_0_159), .Q(QuotientVar[2]), 
      .QN());
   DFF_X1 \QuotientVar_reg[1]  (.D(n_0_116), .CK(n_0_159), .Q(QuotientVar[1]), 
      .QN());
   DFF_X1 \QuotientVar_reg[0]  (.D(n_0_115), .CK(n_0_159), .Q(QuotientVar[0]), 
      .QN());
   DFF_X1 \Divisor2_reg[28]  (.D(n_0_114), .CK(n_0_159), .Q(n_0_35), .QN());
   DFF_X1 \Divisor2_reg[27]  (.D(n_0_113), .CK(n_0_159), .Q(n_0_36), .QN());
   DFF_X1 \Divisor2_reg[26]  (.D(n_0_112), .CK(n_0_159), .Q(n_0_37), .QN());
   DFF_X1 \Divisor2_reg[25]  (.D(n_0_111), .CK(n_0_159), .Q(n_0_38), .QN());
   DFF_X1 \Divisor2_reg[24]  (.D(n_0_110), .CK(n_0_159), .Q(n_0_39), .QN());
   DFF_X1 \Divisor2_reg[23]  (.D(n_0_109), .CK(n_0_159), .Q(n_0_40), .QN());
   DFF_X1 \Divisor2_reg[22]  (.D(n_0_108), .CK(n_0_159), .Q(n_0_41), .QN());
   DFF_X1 \Divisor2_reg[21]  (.D(n_0_107), .CK(n_0_159), .Q(n_0_42), .QN());
   DFF_X1 \Divisor2_reg[20]  (.D(n_0_106), .CK(n_0_159), .Q(n_0_43), .QN());
   DFF_X1 \Divisor2_reg[19]  (.D(n_0_105), .CK(n_0_159), .Q(n_0_44), .QN());
   DFF_X1 \Divisor2_reg[18]  (.D(n_0_104), .CK(n_0_159), .Q(n_0_45), .QN());
   DFF_X1 \Divisor2_reg[17]  (.D(n_0_103), .CK(n_0_159), .Q(n_0_46), .QN());
   DFF_X1 \Divisor2_reg[16]  (.D(n_0_102), .CK(n_0_159), .Q(n_0_47), .QN());
   DFF_X1 \Divisor2_reg[15]  (.D(n_0_101), .CK(n_0_159), .Q(n_0_48), .QN());
   DFF_X1 \Divisor2_reg[14]  (.D(n_0_100), .CK(n_0_159), .Q(n_0_49), .QN());
   DFF_X1 \Divisor2_reg[13]  (.D(n_0_99), .CK(n_0_159), .Q(n_0_50), .QN());
   DFF_X1 \Divisor2_reg[12]  (.D(n_0_98), .CK(n_0_159), .Q(n_0_51), .QN());
   DFF_X1 \Divisor2_reg[11]  (.D(n_0_97), .CK(n_0_159), .Q(n_0_52), .QN());
   DFF_X1 \Divisor2_reg[10]  (.D(n_0_96), .CK(n_0_159), .Q(n_0_53), .QN());
   DFF_X1 \Divisor2_reg[9]  (.D(n_0_95), .CK(n_0_159), .Q(n_0_54), .QN());
   DFF_X1 \Divisor2_reg[8]  (.D(n_0_94), .CK(n_0_159), .Q(n_0_55), .QN());
   DFF_X1 \Divisor2_reg[7]  (.D(n_0_93), .CK(n_0_159), .Q(n_0_56), .QN());
   DFF_X1 \Divisor2_reg[6]  (.D(n_0_92), .CK(n_0_159), .Q(n_0_57), .QN());
   DFF_X1 \Divisor2_reg[5]  (.D(n_0_91), .CK(n_0_159), .Q(n_0_58), .QN());
   DFF_X1 \Divisor2_reg[4]  (.D(n_0_90), .CK(n_0_159), .Q(n_0_59), .QN());
   DFF_X1 \Divisor2_reg[3]  (.D(n_0_89), .CK(n_0_159), .Q(n_0_60), .QN());
   DFF_X1 \Divisor2_reg[2]  (.D(n_0_88), .CK(n_0_159), .Q(n_0_61), .QN());
   DFF_X1 \Divisor2_reg[1]  (.D(n_0_87), .CK(n_0_159), .Q(n_0_62), .QN());
   DFF_X1 \Divisor2_reg[0]  (.D(n_0_86), .CK(n_0_159), .Q(n_0_63), .QN());
   DFF_X1 \Dividend2_reg[14]  (.D(n_0_84), .CK(n_0_0), .Q(Dividend2[14]), .QN());
   DFF_X1 \Dividend2_reg[13]  (.D(n_0_83), .CK(n_0_0), .Q(Dividend2[13]), .QN());
   DFF_X1 \Dividend2_reg[12]  (.D(n_0_82), .CK(n_0_0), .Q(Dividend2[12]), .QN());
   DFF_X1 \Dividend2_reg[11]  (.D(n_0_81), .CK(n_0_0), .Q(Dividend2[11]), .QN());
   DFF_X1 \Dividend2_reg[10]  (.D(n_0_80), .CK(n_0_0), .Q(Dividend2[10]), .QN());
   DFF_X1 \Dividend2_reg[9]  (.D(n_0_79), .CK(n_0_0), .Q(Dividend2[9]), .QN());
   DFF_X1 \Dividend2_reg[8]  (.D(n_0_78), .CK(n_0_0), .Q(Dividend2[8]), .QN());
   DFF_X1 \Dividend2_reg[7]  (.D(n_0_77), .CK(n_0_0), .Q(Dividend2[7]), .QN());
   DFF_X1 \Dividend2_reg[6]  (.D(n_0_76), .CK(n_0_0), .Q(Dividend2[6]), .QN());
   DFF_X1 \Dividend2_reg[5]  (.D(n_0_75), .CK(n_0_0), .Q(Dividend2[5]), .QN());
   DFF_X1 \Dividend2_reg[4]  (.D(n_0_74), .CK(n_0_0), .Q(Dividend2[4]), .QN());
   DFF_X1 \Dividend2_reg[3]  (.D(n_0_73), .CK(n_0_0), .Q(Dividend2[3]), .QN());
   DFF_X1 \Dividend2_reg[2]  (.D(n_0_72), .CK(n_0_0), .Q(Dividend2[2]), .QN());
   DFF_X1 \Dividend2_reg[1]  (.D(n_0_71), .CK(n_0_0), .Q(Dividend2[1]), .QN());
   CLKGATETST_X1 clk_gate_Dividend2_reg__14 (.CK(clk), .E(n_0_68), .SE(1'b0), 
      .GCK(n_0_0));
   DFF_X1 \Dividend2_reg[0]  (.D(n_0_70), .CK(n_0_0), .Q(Dividend2[0]), .QN());
   DFF_X1 \Dividend2_reg[15]  (.D(n_0_64), .CK(clk), .Q(Dividend2[15]), .QN());
   MUX2_X1 \Dividend2_reg[15]_enable_mux_0  (.A(Dividend2[15]), .B(n_0_85), 
      .S(n_0_69), .Z(n_0_64));
   DFF_X1 FIRST_ONE_reg (.D(n_0_65), .CK(clk), .Q(FIRST_ONE), .QN());
   MUX2_X1 FIRST_ONE_reg_enable_mux_0 (.A(FIRST_ONE), .B(n_0_67), .S(n_0_66), 
      .Z(n_0_65));
   CLKGATETST_X1 clk_gate_Done_bit_reg (.CK(clk), .E(n_0_130), .SE(1'b0), 
      .GCK(n_0_159));
   CLKGATETST_X1 clk_gate_add1_reg (.CK(clk), .E(n_0_182), .SE(1'b0), .GCK(
      n_0_142));
   HA_X1 i_0_0_0 (.A(n_0_0_13), .B(n_0_0_14), .CO(n_0_0_19), .S());
   FA_X1 i_0_0_1 (.A(n_0_0_15), .B(n_0_0_16), .CI(n_0_0_19), .CO(n_0_0_20), 
      .S());
   HA_X1 i_0_0_2 (.A(n_0_0_9), .B(n_0_0_17), .CO(n_0_0_0), .S());
   HA_X1 i_0_0_3 (.A(n_0_0_6), .B(n_0_0_0), .CO(n_0_0_1), .S());
   OAI21_X1 i_0_0_4 (.A(n_0_0_2), .B1(n_0_0_283), .B2(n_0_0_306), .ZN(n_0_0_16));
   AOI21_X1 i_0_0_5 (.A(n_0_0_279), .B1(n_0_0_283), .B2(n_0_0_306), .ZN(n_0_0_2));
   XNOR2_X1 i_0_0_6 (.A(n_0_0_5), .B(n_0_0_3), .ZN(n_0_0_14));
   OR2_X1 i_0_0_7 (.A1(n_0_0_5), .A2(n_0_0_3), .ZN(n_0_0_15));
   XNOR2_X1 i_0_0_8 (.A(n_0_0_306), .B(n_0_0_279), .ZN(n_0_0_3));
   OAI211_X1 i_0_0_9 (.A(n_0_0_5), .B(n_0_0_4), .C1(n_0_0_12), .C2(n_0_0_8), 
      .ZN(n_0_0_13));
   AOI22_X1 i_0_0_10 (.A1(n_0_0_9), .A2(n_0_0_290), .B1(n_0_0_294), .B2(n_0_0_6), 
      .ZN(n_0_0_4));
   OR2_X1 i_0_0_11 (.A1(n_0_0_6), .A2(n_0_0_294), .ZN(n_0_0_5));
   OR3_X1 i_0_0_12 (.A1(Divisor[14]), .A2(n_0_0_7), .A3(n_0_0_280), .ZN(n_0_0_6));
   AOI21_X1 i_0_0_13 (.A(n_0_0_281), .B1(n_0_0_285), .B2(n_0_0_287), .ZN(n_0_0_7));
   OAI211_X1 i_0_0_14 (.A(n_0_0_301), .B(n_0_0_298), .C1(n_0_0_9), .C2(n_0_0_290), 
      .ZN(n_0_0_8));
   OAI221_X1 i_0_0_15 (.A(n_0_0_337), .B1(n_0_0_282), .B2(n_0_0_280), .C1(
      n_0_0_10), .C2(n_0_0_279), .ZN(n_0_0_9));
   NOR3_X1 i_0_0_16 (.A1(Divisor[7]), .A2(Divisor[6]), .A3(n_0_0_11), .ZN(
      n_0_0_10));
   NOR3_X1 i_0_0_17 (.A1(Divisor[5]), .A2(Divisor[4]), .A3(n_0_0_288), .ZN(
      n_0_0_11));
   INV_X1 i_0_0_18 (.A(n_0_0_17), .ZN(n_0_0_12));
   NOR2_X1 i_0_0_19 (.A1(Divisor[14]), .A2(n_0_0_18), .ZN(n_0_0_17));
   NOR2_X1 i_0_0_20 (.A1(Divisor[13]), .A2(n_0_0_21), .ZN(n_0_0_18));
   NOR2_X1 i_0_0_21 (.A1(Divisor[12]), .A2(n_0_0_22), .ZN(n_0_0_21));
   AOI21_X1 i_0_0_22 (.A(Divisor[11]), .B1(n_0_0_336), .B2(n_0_0_23), .ZN(
      n_0_0_22));
   OAI21_X1 i_0_0_23 (.A(n_0_0_335), .B1(Divisor[8]), .B2(n_0_0_24), .ZN(
      n_0_0_23));
   AOI21_X1 i_0_0_24 (.A(Divisor[7]), .B1(n_0_0_333), .B2(n_0_0_25), .ZN(
      n_0_0_24));
   OAI21_X1 i_0_0_25 (.A(n_0_0_332), .B1(Divisor[4]), .B2(n_0_0_26), .ZN(
      n_0_0_25));
   AOI21_X1 i_0_0_26 (.A(Divisor[3]), .B1(n_0_0_331), .B2(Divisor[1]), .ZN(
      n_0_0_26));
   AOI21_X1 i_0_0_27 (.A(n_0_0_27), .B1(n_0_0_275), .B2(n_0_0_276), .ZN(n_0_66));
   NOR3_X1 i_0_0_28 (.A1(FIRST_ONE), .A2(n_0_0_172), .A3(n_0_0_263), .ZN(
      n_0_0_27));
   OAI21_X1 i_0_0_29 (.A(n_0_0_275), .B1(n_0_0_102), .B2(Dividend[15]), .ZN(
      n_0_69));
   NAND2_X1 i_0_0_30 (.A1(n_0_0_102), .A2(n_0_0_275), .ZN(n_0_68));
   OAI21_X1 i_0_0_31 (.A(n_0_0_108), .B1(n_0_0_233), .B2(n_0_0_263), .ZN(n_0_70));
   OAI22_X1 i_0_0_32 (.A1(n_0_0_273), .A2(n_0_0_28), .B1(n_0_0_235), .B2(
      n_0_0_263), .ZN(n_0_71));
   XNOR2_X1 i_0_0_33 (.A(n_0_0_339), .B(n_0_0_29), .ZN(n_0_0_28));
   NAND2_X1 i_0_0_34 (.A1(Dividend[15]), .A2(Dividend[0]), .ZN(n_0_0_29));
   OAI22_X1 i_0_0_35 (.A1(n_0_0_273), .A2(n_0_0_30), .B1(n_0_0_230), .B2(
      n_0_0_263), .ZN(n_0_72));
   XNOR2_X1 i_0_0_36 (.A(n_0_0_340), .B(n_0_0_33), .ZN(n_0_0_30));
   OAI22_X1 i_0_0_37 (.A1(n_0_0_273), .A2(n_0_0_31), .B1(n_0_0_227), .B2(
      n_0_0_263), .ZN(n_0_73));
   XNOR2_X1 i_0_0_38 (.A(Dividend[3]), .B(n_0_0_32), .ZN(n_0_0_31));
   AOI21_X1 i_0_0_39 (.A(n_0_0_353), .B1(n_0_0_340), .B2(n_0_0_33), .ZN(n_0_0_32));
   OAI21_X1 i_0_0_40 (.A(Dividend[15]), .B1(Dividend[1]), .B2(Dividend[0]), 
      .ZN(n_0_0_33));
   OAI22_X1 i_0_0_41 (.A1(n_0_0_273), .A2(n_0_0_34), .B1(n_0_0_223), .B2(
      n_0_0_263), .ZN(n_0_74));
   XNOR2_X1 i_0_0_42 (.A(n_0_0_342), .B(n_0_0_43), .ZN(n_0_0_34));
   OAI22_X1 i_0_0_43 (.A1(n_0_0_40), .A2(n_0_0_35), .B1(n_0_0_263), .B2(
      n_0_0_238), .ZN(n_0_75));
   OAI21_X1 i_0_0_44 (.A(n_0_0_274), .B1(n_0_0_42), .B2(n_0_0_343), .ZN(n_0_0_35));
   OAI22_X1 i_0_0_45 (.A1(n_0_0_273), .A2(n_0_0_36), .B1(n_0_0_218), .B2(
      n_0_0_263), .ZN(n_0_76));
   XNOR2_X1 i_0_0_46 (.A(n_0_0_344), .B(n_0_0_39), .ZN(n_0_0_36));
   OAI22_X1 i_0_0_47 (.A1(n_0_0_273), .A2(n_0_0_37), .B1(n_0_0_215), .B2(
      n_0_0_263), .ZN(n_0_77));
   XNOR2_X1 i_0_0_48 (.A(n_0_0_345), .B(n_0_0_38), .ZN(n_0_0_37));
   OAI21_X1 i_0_0_49 (.A(Dividend[15]), .B1(n_0_0_41), .B2(Dividend[6]), 
      .ZN(n_0_0_38));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_41), .A2(Dividend[15]), .ZN(n_0_0_39));
   INV_X1 i_0_0_51 (.A(n_0_0_41), .ZN(n_0_0_40));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_343), .A2(n_0_0_42), .ZN(n_0_0_41));
   OAI21_X1 i_0_0_53 (.A(Dividend[15]), .B1(n_0_0_271), .B2(Dividend[4]), 
      .ZN(n_0_0_42));
   NAND2_X1 i_0_0_54 (.A1(n_0_0_271), .A2(Dividend[15]), .ZN(n_0_0_43));
   OAI22_X1 i_0_0_55 (.A1(n_0_0_273), .A2(n_0_0_44), .B1(n_0_0_212), .B2(
      n_0_0_263), .ZN(n_0_78));
   XNOR2_X1 i_0_0_56 (.A(n_0_0_346), .B(n_0_0_58), .ZN(n_0_0_44));
   OAI21_X1 i_0_0_57 (.A(n_0_0_45), .B1(n_0_0_208), .B2(n_0_0_263), .ZN(n_0_79));
   NAND3_X1 i_0_0_58 (.A1(n_0_0_51), .A2(n_0_0_46), .A3(n_0_0_274), .ZN(n_0_0_45));
   OAI211_X1 i_0_0_59 (.A(Dividend[15]), .B(Dividend[9]), .C1(n_0_0_269), 
      .C2(Dividend[8]), .ZN(n_0_0_46));
   OAI22_X1 i_0_0_60 (.A1(n_0_0_273), .A2(n_0_0_47), .B1(n_0_0_205), .B2(
      n_0_0_263), .ZN(n_0_80));
   XNOR2_X1 i_0_0_61 (.A(n_0_0_348), .B(n_0_0_50), .ZN(n_0_0_47));
   OAI22_X1 i_0_0_62 (.A1(n_0_0_273), .A2(n_0_0_48), .B1(n_0_0_202), .B2(
      n_0_0_263), .ZN(n_0_81));
   XNOR2_X1 i_0_0_63 (.A(n_0_0_349), .B(n_0_0_49), .ZN(n_0_0_48));
   OAI21_X1 i_0_0_64 (.A(Dividend[15]), .B1(n_0_0_51), .B2(Dividend[10]), 
      .ZN(n_0_0_49));
   NAND2_X1 i_0_0_65 (.A1(n_0_0_51), .A2(Dividend[15]), .ZN(n_0_0_50));
   OAI211_X1 i_0_0_66 (.A(n_0_0_347), .B(n_0_0_58), .C1(n_0_0_346), .C2(
      n_0_0_353), .ZN(n_0_0_51));
   OAI22_X1 i_0_0_67 (.A1(n_0_0_273), .A2(n_0_0_52), .B1(n_0_0_198), .B2(
      n_0_0_263), .ZN(n_0_82));
   XNOR2_X1 i_0_0_68 (.A(Dividend[12]), .B(n_0_0_57), .ZN(n_0_0_52));
   OAI22_X1 i_0_0_69 (.A1(n_0_0_273), .A2(n_0_0_53), .B1(n_0_0_195), .B2(
      n_0_0_263), .ZN(n_0_83));
   XNOR2_X1 i_0_0_70 (.A(n_0_0_351), .B(n_0_0_54), .ZN(n_0_0_53));
   AOI21_X1 i_0_0_71 (.A(n_0_0_57), .B1(Dividend[12]), .B2(Dividend[15]), 
      .ZN(n_0_0_54));
   OAI22_X1 i_0_0_72 (.A1(n_0_0_273), .A2(n_0_0_55), .B1(n_0_0_192), .B2(
      n_0_0_263), .ZN(n_0_84));
   XNOR2_X1 i_0_0_73 (.A(n_0_0_352), .B(n_0_0_56), .ZN(n_0_0_55));
   AOI21_X1 i_0_0_74 (.A(n_0_0_57), .B1(n_0_0_307), .B2(Dividend[15]), .ZN(
      n_0_0_56));
   OAI21_X1 i_0_0_75 (.A(n_0_0_58), .B1(n_0_0_308), .B2(n_0_0_353), .ZN(n_0_0_57));
   NAND2_X1 i_0_0_76 (.A1(n_0_0_269), .A2(Dividend[15]), .ZN(n_0_0_58));
   OAI22_X1 i_0_0_77 (.A1(n_0_0_353), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_188), .ZN(n_0_85));
   AND2_X1 i_0_0_78 (.A1(n_0_62), .A2(n_0_0_356), .ZN(n_0_86));
   AND2_X1 i_0_0_79 (.A1(n_0_61), .A2(n_0_0_356), .ZN(n_0_87));
   AND2_X1 i_0_0_80 (.A1(n_0_60), .A2(n_0_0_356), .ZN(n_0_88));
   AND2_X1 i_0_0_81 (.A1(n_0_59), .A2(n_0_0_356), .ZN(n_0_89));
   AND2_X1 i_0_0_82 (.A1(n_0_58), .A2(n_0_0_356), .ZN(n_0_90));
   AND2_X1 i_0_0_83 (.A1(n_0_57), .A2(n_0_0_356), .ZN(n_0_91));
   AND2_X1 i_0_0_84 (.A1(n_0_56), .A2(n_0_0_356), .ZN(n_0_92));
   AND2_X1 i_0_0_85 (.A1(n_0_55), .A2(n_0_0_356), .ZN(n_0_93));
   AND2_X1 i_0_0_86 (.A1(n_0_54), .A2(n_0_0_356), .ZN(n_0_94));
   AND2_X1 i_0_0_87 (.A1(n_0_53), .A2(n_0_0_356), .ZN(n_0_95));
   AND2_X1 i_0_0_88 (.A1(n_0_52), .A2(n_0_0_356), .ZN(n_0_96));
   AND2_X1 i_0_0_89 (.A1(n_0_51), .A2(n_0_0_356), .ZN(n_0_97));
   AND2_X1 i_0_0_90 (.A1(n_0_50), .A2(n_0_0_356), .ZN(n_0_98));
   AND2_X1 i_0_0_91 (.A1(n_0_49), .A2(n_0_0_356), .ZN(n_0_99));
   OAI21_X1 i_0_0_92 (.A(n_0_0_59), .B1(n_0_0_101), .B2(n_0_0_329), .ZN(n_0_100));
   NAND2_X1 i_0_0_93 (.A1(n_0_48), .A2(n_0_0_356), .ZN(n_0_0_59));
   OAI21_X1 i_0_0_94 (.A(n_0_0_62), .B1(n_0_0_101), .B2(n_0_0_60), .ZN(n_0_101));
   XNOR2_X1 i_0_0_95 (.A(n_0_0_330), .B(n_0_0_61), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_96 (.A1(Divisor[15]), .A2(Divisor[0]), .ZN(n_0_0_61));
   NAND2_X1 i_0_0_97 (.A1(n_0_47), .A2(n_0_0_356), .ZN(n_0_0_62));
   OAI21_X1 i_0_0_98 (.A(n_0_0_64), .B1(n_0_0_63), .B2(n_0_0_101), .ZN(n_0_102));
   XNOR2_X1 i_0_0_99 (.A(n_0_0_331), .B(n_0_0_68), .ZN(n_0_0_63));
   NAND2_X1 i_0_0_100 (.A1(n_0_46), .A2(n_0_0_356), .ZN(n_0_0_64));
   OAI21_X1 i_0_0_101 (.A(n_0_0_69), .B1(n_0_0_101), .B2(n_0_0_65), .ZN(n_0_103));
   XOR2_X1 i_0_0_102 (.A(Divisor[3]), .B(n_0_0_66), .Z(n_0_0_65));
   OAI21_X1 i_0_0_103 (.A(Divisor[15]), .B1(Divisor[2]), .B2(n_0_0_67), .ZN(
      n_0_0_66));
   INV_X1 i_0_0_104 (.A(n_0_0_68), .ZN(n_0_0_67));
   OAI21_X1 i_0_0_105 (.A(Divisor[15]), .B1(Divisor[1]), .B2(Divisor[0]), 
      .ZN(n_0_0_68));
   NAND2_X1 i_0_0_106 (.A1(n_0_45), .A2(n_0_0_356), .ZN(n_0_0_69));
   OAI21_X1 i_0_0_107 (.A(n_0_0_71), .B1(n_0_0_70), .B2(n_0_0_101), .ZN(n_0_104));
   XOR2_X1 i_0_0_108 (.A(Divisor[4]), .B(n_0_0_74), .Z(n_0_0_70));
   NAND2_X1 i_0_0_109 (.A1(n_0_44), .A2(n_0_0_356), .ZN(n_0_0_71));
   OAI21_X1 i_0_0_110 (.A(n_0_0_75), .B1(n_0_0_101), .B2(n_0_0_72), .ZN(n_0_105));
   XNOR2_X1 i_0_0_111 (.A(n_0_0_332), .B(n_0_0_73), .ZN(n_0_0_72));
   OAI21_X1 i_0_0_112 (.A(Divisor[15]), .B1(n_0_0_287), .B2(Divisor[4]), 
      .ZN(n_0_0_73));
   NAND2_X1 i_0_0_113 (.A1(n_0_0_287), .A2(Divisor[15]), .ZN(n_0_0_74));
   NAND2_X1 i_0_0_114 (.A1(n_0_43), .A2(n_0_0_356), .ZN(n_0_0_75));
   OAI21_X1 i_0_0_115 (.A(n_0_0_78), .B1(n_0_0_101), .B2(n_0_0_76), .ZN(n_0_106));
   XNOR2_X1 i_0_0_116 (.A(n_0_0_333), .B(n_0_0_77), .ZN(n_0_0_76));
   NAND2_X1 i_0_0_117 (.A1(n_0_0_286), .A2(Divisor[15]), .ZN(n_0_0_77));
   NAND2_X1 i_0_0_118 (.A1(n_0_42), .A2(n_0_0_356), .ZN(n_0_0_78));
   OAI21_X1 i_0_0_119 (.A(n_0_0_81), .B1(n_0_0_79), .B2(n_0_0_101), .ZN(n_0_107));
   XOR2_X1 i_0_0_120 (.A(Divisor[7]), .B(n_0_0_80), .Z(n_0_0_79));
   NAND2_X1 i_0_0_121 (.A1(n_0_0_284), .A2(Divisor[15]), .ZN(n_0_0_80));
   NAND2_X1 i_0_0_122 (.A1(n_0_41), .A2(n_0_0_356), .ZN(n_0_0_81));
   OAI21_X1 i_0_0_123 (.A(n_0_0_83), .B1(n_0_0_82), .B2(n_0_0_101), .ZN(n_0_108));
   XNOR2_X1 i_0_0_124 (.A(n_0_0_334), .B(n_0_0_93), .ZN(n_0_0_82));
   NAND2_X1 i_0_0_125 (.A1(n_0_40), .A2(n_0_0_356), .ZN(n_0_0_83));
   OAI21_X1 i_0_0_126 (.A(n_0_0_85), .B1(n_0_0_84), .B2(n_0_0_101), .ZN(n_0_109));
   XNOR2_X1 i_0_0_127 (.A(n_0_0_335), .B(n_0_0_92), .ZN(n_0_0_84));
   NAND2_X1 i_0_0_128 (.A1(n_0_39), .A2(n_0_0_356), .ZN(n_0_0_85));
   OAI21_X1 i_0_0_129 (.A(n_0_0_87), .B1(n_0_0_86), .B2(n_0_0_101), .ZN(n_0_110));
   XNOR2_X1 i_0_0_130 (.A(n_0_0_336), .B(n_0_0_90), .ZN(n_0_0_86));
   NAND2_X1 i_0_0_131 (.A1(n_0_38), .A2(n_0_0_356), .ZN(n_0_0_87));
   OAI21_X1 i_0_0_132 (.A(n_0_0_94), .B1(n_0_0_88), .B2(n_0_0_101), .ZN(n_0_111));
   XOR2_X1 i_0_0_133 (.A(Divisor[11]), .B(n_0_0_89), .Z(n_0_0_88));
   OAI21_X1 i_0_0_134 (.A(Divisor[15]), .B1(n_0_0_91), .B2(Divisor[10]), 
      .ZN(n_0_0_89));
   NAND2_X1 i_0_0_135 (.A1(n_0_0_91), .A2(Divisor[15]), .ZN(n_0_0_90));
   NAND2_X1 i_0_0_136 (.A1(n_0_0_335), .A2(n_0_0_92), .ZN(n_0_0_91));
   OAI21_X1 i_0_0_137 (.A(Divisor[15]), .B1(n_0_0_283), .B2(Divisor[8]), 
      .ZN(n_0_0_92));
   NAND2_X1 i_0_0_138 (.A1(n_0_0_283), .A2(Divisor[15]), .ZN(n_0_0_93));
   NAND2_X1 i_0_0_139 (.A1(n_0_37), .A2(n_0_0_356), .ZN(n_0_0_94));
   OAI21_X1 i_0_0_140 (.A(n_0_0_96), .B1(n_0_0_95), .B2(n_0_0_101), .ZN(n_0_112));
   XOR2_X1 i_0_0_141 (.A(Divisor[12]), .B(n_0_0_104), .Z(n_0_0_95));
   NAND2_X1 i_0_0_142 (.A1(n_0_36), .A2(n_0_0_356), .ZN(n_0_0_96));
   OAI21_X1 i_0_0_143 (.A(n_0_0_99), .B1(n_0_0_97), .B2(n_0_0_101), .ZN(n_0_113));
   XOR2_X1 i_0_0_144 (.A(Divisor[13]), .B(n_0_0_98), .Z(n_0_0_97));
   OAI21_X1 i_0_0_145 (.A(Divisor[15]), .B1(n_0_0_105), .B2(Divisor[12]), 
      .ZN(n_0_0_98));
   NAND2_X1 i_0_0_146 (.A1(n_0_35), .A2(n_0_0_356), .ZN(n_0_0_99));
   NOR2_X1 i_0_0_147 (.A1(n_0_0_101), .A2(n_0_0_100), .ZN(n_0_114));
   XNOR2_X1 i_0_0_148 (.A(n_0_0_337), .B(n_0_0_103), .ZN(n_0_0_100));
   NAND2_X1 i_0_0_149 (.A1(n_0_0_274), .A2(n_0_0_266), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_150 (.A1(Start), .A2(n_0_0_266), .ZN(n_0_0_102));
   OAI21_X1 i_0_0_151 (.A(Divisor[15]), .B1(n_0_0_280), .B2(n_0_0_105), .ZN(
      n_0_0_103));
   NAND2_X1 i_0_0_152 (.A1(n_0_0_105), .A2(Divisor[15]), .ZN(n_0_0_104));
   OR2_X1 i_0_0_153 (.A1(n_0_0_283), .A2(n_0_0_281), .ZN(n_0_0_105));
   OAI22_X1 i_0_0_154 (.A1(n_0_0_145), .A2(n_0_0_263), .B1(n_0_0_338), .B2(
      n_0_0_106), .ZN(n_0_115));
   OAI22_X1 i_0_0_155 (.A1(n_0_0_146), .A2(n_0_0_263), .B1(n_0_0_339), .B2(
      n_0_0_106), .ZN(n_0_116));
   OAI22_X1 i_0_0_156 (.A1(n_0_0_147), .A2(n_0_0_263), .B1(n_0_0_340), .B2(
      n_0_0_106), .ZN(n_0_117));
   OAI22_X1 i_0_0_157 (.A1(n_0_0_148), .A2(n_0_0_263), .B1(n_0_0_341), .B2(
      n_0_0_106), .ZN(n_0_118));
   OAI22_X1 i_0_0_158 (.A1(n_0_0_150), .A2(n_0_0_263), .B1(n_0_0_342), .B2(
      n_0_0_106), .ZN(n_0_119));
   OAI22_X1 i_0_0_159 (.A1(n_0_0_151), .A2(n_0_0_263), .B1(n_0_0_343), .B2(
      n_0_0_106), .ZN(n_0_120));
   OAI22_X1 i_0_0_160 (.A1(n_0_0_152), .A2(n_0_0_263), .B1(n_0_0_344), .B2(
      n_0_0_106), .ZN(n_0_121));
   OAI22_X1 i_0_0_161 (.A1(n_0_0_153), .A2(n_0_0_263), .B1(n_0_0_345), .B2(
      n_0_0_106), .ZN(n_0_122));
   OAI22_X1 i_0_0_162 (.A1(n_0_0_156), .A2(n_0_0_263), .B1(n_0_0_346), .B2(
      n_0_0_106), .ZN(n_0_123));
   OAI22_X1 i_0_0_163 (.A1(n_0_0_157), .A2(n_0_0_263), .B1(n_0_0_347), .B2(
      n_0_0_106), .ZN(n_0_124));
   OAI22_X1 i_0_0_164 (.A1(n_0_0_158), .A2(n_0_0_263), .B1(n_0_0_348), .B2(
      n_0_0_106), .ZN(n_0_125));
   OAI22_X1 i_0_0_165 (.A1(n_0_0_162), .A2(n_0_0_263), .B1(n_0_0_349), .B2(
      n_0_0_106), .ZN(n_0_126));
   OAI22_X1 i_0_0_166 (.A1(n_0_0_161), .A2(n_0_0_263), .B1(n_0_0_350), .B2(
      n_0_0_106), .ZN(n_0_127));
   OAI22_X1 i_0_0_167 (.A1(n_0_0_164), .A2(n_0_0_263), .B1(n_0_0_351), .B2(
      n_0_0_106), .ZN(n_0_128));
   OAI22_X1 i_0_0_168 (.A1(n_0_0_143), .A2(n_0_0_263), .B1(n_0_0_352), .B2(
      n_0_0_106), .ZN(n_0_129));
   OR2_X1 i_0_0_169 (.A1(n_0_0_242), .A2(rst), .ZN(n_0_0_106));
   OAI21_X1 i_0_0_170 (.A(n_0_0_272), .B1(n_0_2), .B2(Index[0]), .ZN(n_0_131));
   AND2_X1 i_0_0_171 (.A1(n_0_3), .A2(n_0_0_356), .ZN(n_0_132));
   OAI21_X1 i_0_0_172 (.A(n_0_0_272), .B1(n_0_0_310), .B2(n_0_2), .ZN(n_0_133));
   AND2_X1 i_0_0_173 (.A1(n_0_5), .A2(n_0_0_356), .ZN(n_0_134));
   OAI21_X1 i_0_0_174 (.A(n_0_0_272), .B1(n_0_0_311), .B2(n_0_2), .ZN(n_0_135));
   NAND2_X1 i_0_0_175 (.A1(n_0_0_275), .A2(n_0_0_276), .ZN(n_0_130));
   AND2_X1 i_0_0_176 (.A1(n_0_7), .A2(n_0_0_356), .ZN(n_0_136));
   AND2_X1 i_0_0_177 (.A1(n_0_8), .A2(n_0_0_356), .ZN(n_0_137));
   AND2_X1 i_0_0_178 (.A1(n_0_9), .A2(n_0_0_356), .ZN(n_0_138));
   AND2_X1 i_0_0_179 (.A1(n_0_10), .A2(n_0_0_356), .ZN(n_0_139));
   AND2_X1 i_0_0_180 (.A1(n_0_11), .A2(n_0_0_356), .ZN(n_0_140));
   AND2_X1 i_0_0_181 (.A1(n_0_12), .A2(n_0_0_356), .ZN(n_0_141));
   AND2_X1 i_0_0_182 (.A1(n_0_13), .A2(n_0_0_356), .ZN(n_0_143));
   AND2_X1 i_0_0_183 (.A1(n_0_14), .A2(n_0_0_356), .ZN(n_0_144));
   AND2_X1 i_0_0_184 (.A1(n_0_15), .A2(n_0_0_356), .ZN(n_0_145));
   AND2_X1 i_0_0_185 (.A1(n_0_16), .A2(n_0_0_356), .ZN(n_0_146));
   AND2_X1 i_0_0_186 (.A1(n_0_17), .A2(n_0_0_356), .ZN(n_0_147));
   AND2_X1 i_0_0_187 (.A1(n_0_18), .A2(n_0_0_356), .ZN(n_0_148));
   AND2_X1 i_0_0_188 (.A1(n_0_19), .A2(n_0_0_356), .ZN(n_0_149));
   AND2_X1 i_0_0_189 (.A1(n_0_20), .A2(n_0_0_356), .ZN(n_0_150));
   AND2_X1 i_0_0_190 (.A1(n_0_21), .A2(n_0_0_356), .ZN(n_0_151));
   AND2_X1 i_0_0_191 (.A1(n_0_22), .A2(n_0_0_356), .ZN(n_0_152));
   AND2_X1 i_0_0_192 (.A1(n_0_23), .A2(n_0_0_356), .ZN(n_0_153));
   AND2_X1 i_0_0_193 (.A1(n_0_24), .A2(n_0_0_356), .ZN(n_0_154));
   AND2_X1 i_0_0_194 (.A1(n_0_26), .A2(n_0_0_356), .ZN(n_0_155));
   AND2_X1 i_0_0_195 (.A1(n_0_27), .A2(n_0_0_356), .ZN(n_0_156));
   AND2_X1 i_0_0_196 (.A1(n_0_28), .A2(n_0_0_356), .ZN(n_0_157));
   AND2_X1 i_0_0_197 (.A1(n_0_29), .A2(n_0_0_356), .ZN(n_0_158));
   AND2_X1 i_0_0_198 (.A1(n_0_30), .A2(n_0_0_356), .ZN(n_0_160));
   AND2_X1 i_0_0_199 (.A1(n_0_31), .A2(n_0_0_356), .ZN(n_0_161));
   AND2_X1 i_0_0_200 (.A1(n_0_32), .A2(n_0_0_356), .ZN(n_0_162));
   AND2_X1 i_0_0_201 (.A1(n_0_33), .A2(n_0_0_356), .ZN(n_0_163));
   AND2_X1 i_0_0_202 (.A1(n_0_34), .A2(n_0_0_356), .ZN(n_0_164));
   NAND2_X1 i_0_0_203 (.A1(n_0_0_262), .A2(n_0_0_243), .ZN(n_0_165));
   NOR2_X1 i_0_0_204 (.A1(rst), .A2(n_0_0_233), .ZN(n_0_166));
   NOR2_X1 i_0_0_205 (.A1(rst), .A2(n_0_0_235), .ZN(n_0_167));
   NOR2_X1 i_0_0_206 (.A1(rst), .A2(n_0_0_230), .ZN(n_0_168));
   NOR2_X1 i_0_0_207 (.A1(rst), .A2(n_0_0_227), .ZN(n_0_169));
   NOR2_X1 i_0_0_208 (.A1(rst), .A2(n_0_0_223), .ZN(n_0_170));
   NOR2_X1 i_0_0_209 (.A1(rst), .A2(n_0_0_238), .ZN(n_0_171));
   NOR2_X1 i_0_0_210 (.A1(rst), .A2(n_0_0_218), .ZN(n_0_172));
   NOR2_X1 i_0_0_211 (.A1(rst), .A2(n_0_0_215), .ZN(n_0_173));
   NOR2_X1 i_0_0_212 (.A1(rst), .A2(n_0_0_212), .ZN(n_0_174));
   NOR2_X1 i_0_0_213 (.A1(rst), .A2(n_0_0_208), .ZN(n_0_175));
   NOR2_X1 i_0_0_214 (.A1(rst), .A2(n_0_0_205), .ZN(n_0_176));
   NOR2_X1 i_0_0_215 (.A1(rst), .A2(n_0_0_202), .ZN(n_0_177));
   NOR2_X1 i_0_0_216 (.A1(rst), .A2(n_0_0_198), .ZN(n_0_178));
   NOR2_X1 i_0_0_217 (.A1(rst), .A2(n_0_0_195), .ZN(n_0_179));
   NOR2_X1 i_0_0_218 (.A1(rst), .A2(n_0_0_192), .ZN(n_0_180));
   NOR2_X1 i_0_0_219 (.A1(n_0_0_188), .A2(rst), .ZN(n_0_181));
   INV_X1 i_0_0_220 (.A(n_0_0_107), .ZN(n_0_182));
   NOR2_X1 i_0_0_221 (.A1(rst), .A2(n_0_67), .ZN(n_0_0_107));
   AND3_X1 i_0_0_222 (.A1(n_0_0_187), .A2(n_0_0_174), .A3(n_0_0_356), .ZN(n_0_67));
   NOR2_X1 i_0_0_223 (.A1(n_0_63), .A2(rst), .ZN(n_0_183));
   NOR2_X1 i_0_0_224 (.A1(n_0_62), .A2(rst), .ZN(n_0_184));
   NOR2_X1 i_0_0_225 (.A1(n_0_61), .A2(rst), .ZN(n_0_185));
   NOR2_X1 i_0_0_226 (.A1(n_0_60), .A2(rst), .ZN(n_0_186));
   NOR2_X1 i_0_0_227 (.A1(n_0_59), .A2(rst), .ZN(n_0_187));
   NOR2_X1 i_0_0_228 (.A1(n_0_58), .A2(rst), .ZN(n_0_188));
   NOR2_X1 i_0_0_229 (.A1(n_0_57), .A2(rst), .ZN(n_0_189));
   NOR2_X1 i_0_0_230 (.A1(n_0_56), .A2(rst), .ZN(n_0_190));
   NOR2_X1 i_0_0_231 (.A1(n_0_55), .A2(rst), .ZN(n_0_191));
   NOR2_X1 i_0_0_232 (.A1(n_0_54), .A2(rst), .ZN(n_0_192));
   NOR2_X1 i_0_0_233 (.A1(n_0_53), .A2(rst), .ZN(n_0_193));
   NOR2_X1 i_0_0_234 (.A1(n_0_52), .A2(rst), .ZN(n_0_194));
   NOR2_X1 i_0_0_235 (.A1(n_0_51), .A2(rst), .ZN(n_0_195));
   NOR2_X1 i_0_0_236 (.A1(n_0_50), .A2(rst), .ZN(n_0_196));
   NOR2_X1 i_0_0_237 (.A1(n_0_49), .A2(rst), .ZN(n_0_197));
   NOR2_X1 i_0_0_238 (.A1(n_0_48), .A2(rst), .ZN(n_0_198));
   NAND2_X1 i_0_0_239 (.A1(n_0_0_243), .A2(n_0_0_242), .ZN(n_0_199));
   OAI21_X1 i_0_0_240 (.A(n_0_0_108), .B1(n_0_0_145), .B2(n_0_0_263), .ZN(
      n_0_200));
   NAND2_X1 i_0_0_241 (.A1(Dividend[0]), .A2(n_0_0_274), .ZN(n_0_0_108));
   OAI22_X1 i_0_0_242 (.A1(n_0_0_339), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_109), .ZN(n_0_201));
   XOR2_X1 i_0_0_243 (.A(n_0_0_146), .B(n_0_0_144), .Z(n_0_0_109));
   OAI22_X1 i_0_0_244 (.A1(n_0_0_340), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_110), .ZN(n_0_202));
   XOR2_X1 i_0_0_245 (.A(n_0_0_147), .B(n_0_0_111), .Z(n_0_0_110));
   AOI21_X1 i_0_0_246 (.A(n_0_0_357), .B1(n_0_0_146), .B2(n_0_0_145), .ZN(
      n_0_0_111));
   OAI22_X1 i_0_0_247 (.A1(n_0_0_341), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_112), .ZN(n_0_203));
   XOR2_X1 i_0_0_248 (.A(n_0_0_148), .B(n_0_0_113), .Z(n_0_0_112));
   NOR2_X1 i_0_0_249 (.A1(n_0_0_142), .A2(n_0_0_357), .ZN(n_0_0_113));
   OAI22_X1 i_0_0_250 (.A1(n_0_0_342), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_114), .ZN(n_0_204));
   XNOR2_X1 i_0_0_251 (.A(n_0_0_150), .B(n_0_0_115), .ZN(n_0_0_114));
   NAND2_X1 i_0_0_252 (.A1(n_0_0_141), .A2(n_0_0_166), .ZN(n_0_0_115));
   OAI22_X1 i_0_0_253 (.A1(n_0_0_343), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_116), .ZN(n_0_205));
   XOR2_X1 i_0_0_254 (.A(n_0_0_151), .B(n_0_0_117), .Z(n_0_0_116));
   NOR2_X1 i_0_0_255 (.A1(n_0_0_140), .A2(n_0_0_357), .ZN(n_0_0_117));
   OAI22_X1 i_0_0_256 (.A1(n_0_0_344), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_118), .ZN(n_0_206));
   XOR2_X1 i_0_0_257 (.A(n_0_0_152), .B(n_0_0_119), .Z(n_0_0_118));
   NOR2_X1 i_0_0_258 (.A1(n_0_0_139), .A2(n_0_0_357), .ZN(n_0_0_119));
   OAI22_X1 i_0_0_259 (.A1(n_0_0_345), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_120), .ZN(n_0_207));
   XOR2_X1 i_0_0_260 (.A(n_0_0_153), .B(n_0_0_121), .Z(n_0_0_120));
   AOI21_X1 i_0_0_261 (.A(n_0_0_357), .B1(n_0_0_152), .B2(n_0_0_139), .ZN(
      n_0_0_121));
   OAI22_X1 i_0_0_262 (.A1(n_0_0_346), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_122), .ZN(n_0_208));
   XNOR2_X1 i_0_0_263 (.A(n_0_0_156), .B(n_0_0_123), .ZN(n_0_0_122));
   NAND2_X1 i_0_0_264 (.A1(n_0_0_138), .A2(n_0_0_166), .ZN(n_0_0_123));
   OAI22_X1 i_0_0_265 (.A1(n_0_0_347), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_124), .ZN(n_0_209));
   XOR2_X1 i_0_0_266 (.A(n_0_0_157), .B(n_0_0_125), .Z(n_0_0_124));
   NOR2_X1 i_0_0_267 (.A1(n_0_0_137), .A2(n_0_0_357), .ZN(n_0_0_125));
   OAI22_X1 i_0_0_268 (.A1(n_0_0_348), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_126), .ZN(n_0_210));
   XOR2_X1 i_0_0_269 (.A(n_0_0_158), .B(n_0_0_127), .Z(n_0_0_126));
   AOI21_X1 i_0_0_270 (.A(n_0_0_357), .B1(n_0_0_157), .B2(n_0_0_137), .ZN(
      n_0_0_127));
   OAI22_X1 i_0_0_271 (.A1(n_0_0_349), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_128), .ZN(n_0_211));
   XNOR2_X1 i_0_0_272 (.A(n_0_0_162), .B(n_0_0_135), .ZN(n_0_0_128));
   OAI22_X1 i_0_0_273 (.A1(n_0_0_350), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_129), .ZN(n_0_212));
   XOR2_X1 i_0_0_274 (.A(n_0_0_161), .B(n_0_0_130), .Z(n_0_0_129));
   OAI21_X1 i_0_0_275 (.A(n_0_0_135), .B1(n_0_0_162), .B2(n_0_0_357), .ZN(
      n_0_0_130));
   OAI22_X1 i_0_0_276 (.A1(n_0_0_351), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_131), .ZN(n_0_213));
   XNOR2_X1 i_0_0_277 (.A(n_0_0_164), .B(n_0_0_134), .ZN(n_0_0_131));
   OAI22_X1 i_0_0_278 (.A1(n_0_0_352), .A2(n_0_0_273), .B1(n_0_0_263), .B2(
      n_0_0_132), .ZN(n_0_214));
   XOR2_X1 i_0_0_279 (.A(n_0_0_143), .B(n_0_0_133), .Z(n_0_0_132));
   OAI21_X1 i_0_0_280 (.A(n_0_0_134), .B1(n_0_0_164), .B2(n_0_0_357), .ZN(
      n_0_0_133));
   OAI21_X1 i_0_0_281 (.A(n_0_0_166), .B1(n_0_0_160), .B2(n_0_0_136), .ZN(
      n_0_0_134));
   NAND2_X1 i_0_0_282 (.A1(n_0_0_136), .A2(n_0_0_166), .ZN(n_0_0_135));
   NAND3_X1 i_0_0_283 (.A1(n_0_0_158), .A2(n_0_0_157), .A3(n_0_0_137), .ZN(
      n_0_0_136));
   NOR2_X1 i_0_0_284 (.A1(n_0_0_155), .A2(n_0_0_138), .ZN(n_0_0_137));
   NAND3_X1 i_0_0_285 (.A1(n_0_0_153), .A2(n_0_0_152), .A3(n_0_0_139), .ZN(
      n_0_0_138));
   AND2_X1 i_0_0_286 (.A1(n_0_0_151), .A2(n_0_0_140), .ZN(n_0_0_139));
   AND3_X1 i_0_0_287 (.A1(n_0_0_150), .A2(n_0_0_148), .A3(n_0_0_142), .ZN(
      n_0_0_140));
   NAND2_X1 i_0_0_288 (.A1(n_0_0_148), .A2(n_0_0_142), .ZN(n_0_0_141));
   AND3_X1 i_0_0_289 (.A1(n_0_0_147), .A2(n_0_0_146), .A3(n_0_0_145), .ZN(
      n_0_0_142));
   AOI21_X1 i_0_0_290 (.A(QuotientVar[14]), .B1(n_0_0_169), .B2(n_0_0_159), 
      .ZN(n_0_0_143));
   NOR2_X1 i_0_0_291 (.A1(n_0_0_145), .A2(n_0_0_357), .ZN(n_0_0_144));
   AOI21_X1 i_0_0_292 (.A(QuotientVar[0]), .B1(n_0_0_244), .B2(n_0_0_172), 
      .ZN(n_0_0_145));
   AOI21_X1 i_0_0_293 (.A(QuotientVar[1]), .B1(n_0_0_165), .B2(n_0_0_149), 
      .ZN(n_0_0_146));
   AOI21_X1 i_0_0_294 (.A(QuotientVar[2]), .B1(n_0_0_159), .B2(n_0_0_149), 
      .ZN(n_0_0_147));
   AOI21_X1 i_0_0_295 (.A(QuotientVar[3]), .B1(n_0_0_240), .B2(n_0_0_149), 
      .ZN(n_0_0_148));
   NOR3_X1 i_0_0_296 (.A1(n_0_0_171), .A2(Index[2]), .A3(Index[3]), .ZN(
      n_0_0_149));
   AOI21_X1 i_0_0_297 (.A(QuotientVar[4]), .B1(n_0_0_245), .B2(n_0_0_154), 
      .ZN(n_0_0_150));
   AOI21_X1 i_0_0_298 (.A(QuotientVar[5]), .B1(n_0_0_165), .B2(n_0_0_154), 
      .ZN(n_0_0_151));
   AOI21_X1 i_0_0_299 (.A(QuotientVar[6]), .B1(n_0_0_159), .B2(n_0_0_154), 
      .ZN(n_0_0_152));
   AOI21_X1 i_0_0_300 (.A(QuotientVar[7]), .B1(n_0_0_240), .B2(n_0_0_154), 
      .ZN(n_0_0_153));
   AND3_X1 i_0_0_301 (.A1(n_0_0_170), .A2(n_0_0_355), .A3(Index[2]), .ZN(
      n_0_0_154));
   INV_X1 i_0_0_302 (.A(n_0_0_156), .ZN(n_0_0_155));
   AOI21_X1 i_0_0_303 (.A(QuotientVar[8]), .B1(n_0_0_247), .B2(n_0_0_163), 
      .ZN(n_0_0_156));
   AOI21_X1 i_0_0_304 (.A(QuotientVar[9]), .B1(n_0_0_165), .B2(n_0_0_163), 
      .ZN(n_0_0_157));
   AOI21_X1 i_0_0_305 (.A(QuotientVar[10]), .B1(n_0_0_163), .B2(n_0_0_159), 
      .ZN(n_0_0_158));
   AND2_X1 i_0_0_306 (.A1(n_0_0_354), .A2(Index[1]), .ZN(n_0_0_159));
   NAND2_X1 i_0_0_307 (.A1(n_0_0_162), .A2(n_0_0_161), .ZN(n_0_0_160));
   AOI21_X1 i_0_0_308 (.A(QuotientVar[12]), .B1(n_0_0_247), .B2(n_0_0_169), 
      .ZN(n_0_0_161));
   AOI21_X1 i_0_0_309 (.A(QuotientVar[11]), .B1(n_0_0_240), .B2(n_0_0_163), 
      .ZN(n_0_0_162));
   NOR3_X1 i_0_0_310 (.A1(n_0_0_355), .A2(n_0_0_171), .A3(Index[2]), .ZN(
      n_0_0_163));
   AOI21_X1 i_0_0_311 (.A(QuotientVar[13]), .B1(n_0_0_169), .B2(n_0_0_165), 
      .ZN(n_0_0_164));
   NOR2_X1 i_0_0_312 (.A1(n_0_0_354), .A2(Index[1]), .ZN(n_0_0_165));
   AND2_X1 i_0_0_313 (.A1(QuotientVar[15]), .A2(n_0_0_244), .ZN(n_0_0_166));
   OAI22_X1 i_0_0_314 (.A1(n_0_0_168), .A2(n_0_0_263), .B1(n_0_0_273), .B2(
      n_0_0_167), .ZN(n_0_215));
   XNOR2_X1 i_0_0_315 (.A(Dividend[15]), .B(Divisor[15]), .ZN(n_0_0_167));
   AOI21_X1 i_0_0_316 (.A(QuotientVar[15]), .B1(n_0_0_240), .B2(n_0_0_169), 
      .ZN(n_0_0_168));
   AND3_X1 i_0_0_317 (.A1(Index[3]), .A2(Index[2]), .A3(n_0_0_170), .ZN(
      n_0_0_169));
   INV_X1 i_0_0_318 (.A(n_0_0_171), .ZN(n_0_0_170));
   NAND2_X1 i_0_0_319 (.A1(n_0_0_248), .A2(n_0_0_172), .ZN(n_0_0_171));
   AOI211_X1 i_0_0_320 (.A(n_0_0_176), .B(n_0_0_173), .C1(n_0_0_184), .C2(
      n_0_0_181), .ZN(n_0_0_172));
   NAND2_X1 i_0_0_321 (.A1(n_0_0_187), .A2(n_0_0_175), .ZN(n_0_0_173));
   AOI221_X1 i_0_0_322 (.A(n_0_0_176), .B1(n_0_0_188), .B2(n_0_48), .C1(
      n_0_0_184), .C2(n_0_0_181), .ZN(n_0_0_174));
   NAND2_X1 i_0_0_323 (.A1(n_0_0_188), .A2(n_0_48), .ZN(n_0_0_175));
   NAND4_X1 i_0_0_324 (.A1(n_0_0_180), .A2(n_0_0_179), .A3(n_0_0_178), .A4(
      n_0_0_177), .ZN(n_0_0_176));
   NOR4_X1 i_0_0_325 (.A1(n_0_41), .A2(n_0_42), .A3(n_0_43), .A4(n_0_44), 
      .ZN(n_0_0_177));
   NOR3_X1 i_0_0_326 (.A1(n_0_45), .A2(n_0_46), .A3(n_0_47), .ZN(n_0_0_178));
   NOR2_X1 i_0_0_327 (.A1(n_0_35), .A2(n_0_36), .ZN(n_0_0_179));
   NOR4_X1 i_0_0_328 (.A1(n_0_37), .A2(n_0_38), .A3(n_0_39), .A4(n_0_40), 
      .ZN(n_0_0_180));
   NOR2_X1 i_0_0_329 (.A1(n_0_0_183), .A2(n_0_0_182), .ZN(n_0_0_181));
   NAND4_X1 i_0_0_330 (.A1(n_0_0_212), .A2(n_0_0_208), .A3(n_0_0_205), .A4(
      n_0_0_202), .ZN(n_0_0_182));
   NAND4_X1 i_0_0_331 (.A1(n_0_0_198), .A2(n_0_0_195), .A3(n_0_0_192), .A4(
      n_0_0_188), .ZN(n_0_0_183));
   NOR2_X1 i_0_0_332 (.A1(n_0_0_186), .A2(n_0_0_185), .ZN(n_0_0_184));
   NAND4_X1 i_0_0_333 (.A1(n_0_0_238), .A2(n_0_0_235), .A3(n_0_0_233), .A4(
      n_0_0_230), .ZN(n_0_0_185));
   NAND4_X1 i_0_0_334 (.A1(n_0_0_227), .A2(n_0_0_223), .A3(n_0_0_218), .A4(
      n_0_0_215), .ZN(n_0_0_186));
   OAI221_X1 i_0_0_335 (.A(n_0_0_190), .B1(n_0_0_188), .B2(n_0_48), .C1(n_0_49), 
      .C2(n_0_0_192), .ZN(n_0_0_187));
   OAI21_X1 i_0_0_336 (.A(n_0_0_189), .B1(FIRST_ONE), .B2(Dividend2[15]), 
      .ZN(n_0_0_188));
   NAND2_X1 i_0_0_337 (.A1(n_0_0_327), .A2(FIRST_ONE), .ZN(n_0_0_189));
   OAI21_X1 i_0_0_338 (.A(n_0_0_191), .B1(n_0_0_197), .B2(n_0_0_194), .ZN(
      n_0_0_190));
   AOI22_X1 i_0_0_339 (.A1(n_0_50), .A2(n_0_0_195), .B1(n_0_0_192), .B2(n_0_49), 
      .ZN(n_0_0_191));
   OAI21_X1 i_0_0_340 (.A(n_0_0_193), .B1(FIRST_ONE), .B2(Dividend2[14]), 
      .ZN(n_0_0_192));
   NAND2_X1 i_0_0_341 (.A1(n_0_0_326), .A2(FIRST_ONE), .ZN(n_0_0_193));
   OAI22_X1 i_0_0_342 (.A1(n_0_51), .A2(n_0_0_198), .B1(n_0_0_195), .B2(n_0_50), 
      .ZN(n_0_0_194));
   OAI21_X1 i_0_0_343 (.A(n_0_0_196), .B1(FIRST_ONE), .B2(Dividend2[13]), 
      .ZN(n_0_0_195));
   NAND2_X1 i_0_0_344 (.A1(n_0_0_325), .A2(FIRST_ONE), .ZN(n_0_0_196));
   AOI221_X1 i_0_0_345 (.A(n_0_0_200), .B1(n_0_0_198), .B2(n_0_51), .C1(n_0_52), 
      .C2(n_0_0_202), .ZN(n_0_0_197));
   OAI21_X1 i_0_0_346 (.A(n_0_0_199), .B1(FIRST_ONE), .B2(Dividend2[12]), 
      .ZN(n_0_0_198));
   NAND2_X1 i_0_0_347 (.A1(n_0_0_324), .A2(FIRST_ONE), .ZN(n_0_0_199));
   AOI21_X1 i_0_0_348 (.A(n_0_0_201), .B1(n_0_0_207), .B2(n_0_0_204), .ZN(
      n_0_0_200));
   OAI22_X1 i_0_0_349 (.A1(n_0_53), .A2(n_0_0_205), .B1(n_0_0_202), .B2(n_0_52), 
      .ZN(n_0_0_201));
   OAI21_X1 i_0_0_350 (.A(n_0_0_203), .B1(FIRST_ONE), .B2(Dividend2[11]), 
      .ZN(n_0_0_202));
   NAND2_X1 i_0_0_351 (.A1(n_0_0_323), .A2(FIRST_ONE), .ZN(n_0_0_203));
   AOI22_X1 i_0_0_352 (.A1(n_0_54), .A2(n_0_0_208), .B1(n_0_0_205), .B2(n_0_53), 
      .ZN(n_0_0_204));
   OAI21_X1 i_0_0_353 (.A(n_0_0_206), .B1(FIRST_ONE), .B2(Dividend2[10]), 
      .ZN(n_0_0_205));
   NAND2_X1 i_0_0_354 (.A1(n_0_0_322), .A2(FIRST_ONE), .ZN(n_0_0_206));
   OAI221_X1 i_0_0_355 (.A(n_0_0_210), .B1(n_0_0_208), .B2(n_0_54), .C1(n_0_55), 
      .C2(n_0_0_212), .ZN(n_0_0_207));
   OAI21_X1 i_0_0_356 (.A(n_0_0_209), .B1(FIRST_ONE), .B2(Dividend2[9]), 
      .ZN(n_0_0_208));
   NAND2_X1 i_0_0_357 (.A1(n_0_0_321), .A2(FIRST_ONE), .ZN(n_0_0_209));
   OAI21_X1 i_0_0_358 (.A(n_0_0_211), .B1(n_0_0_217), .B2(n_0_0_214), .ZN(
      n_0_0_210));
   AOI22_X1 i_0_0_359 (.A1(n_0_56), .A2(n_0_0_215), .B1(n_0_0_212), .B2(n_0_55), 
      .ZN(n_0_0_211));
   OAI21_X1 i_0_0_360 (.A(n_0_0_213), .B1(FIRST_ONE), .B2(Dividend2[8]), 
      .ZN(n_0_0_212));
   NAND2_X1 i_0_0_361 (.A1(n_0_0_320), .A2(FIRST_ONE), .ZN(n_0_0_213));
   OAI22_X1 i_0_0_362 (.A1(n_0_57), .A2(n_0_0_218), .B1(n_0_0_215), .B2(n_0_56), 
      .ZN(n_0_0_214));
   OAI21_X1 i_0_0_363 (.A(n_0_0_216), .B1(FIRST_ONE), .B2(Dividend2[7]), 
      .ZN(n_0_0_215));
   NAND2_X1 i_0_0_364 (.A1(n_0_0_319), .A2(FIRST_ONE), .ZN(n_0_0_216));
   AOI21_X1 i_0_0_365 (.A(n_0_0_220), .B1(n_0_0_218), .B2(n_0_57), .ZN(n_0_0_217));
   OAI21_X1 i_0_0_366 (.A(n_0_0_219), .B1(FIRST_ONE), .B2(Dividend2[6]), 
      .ZN(n_0_0_218));
   NAND2_X1 i_0_0_367 (.A1(n_0_0_318), .A2(FIRST_ONE), .ZN(n_0_0_219));
   AOI21_X1 i_0_0_368 (.A(n_0_0_237), .B1(n_0_0_222), .B2(n_0_0_221), .ZN(
      n_0_0_220));
   AOI22_X1 i_0_0_369 (.A1(n_0_58), .A2(n_0_0_238), .B1(n_0_0_223), .B2(n_0_59), 
      .ZN(n_0_0_221));
   OAI221_X1 i_0_0_370 (.A(n_0_0_225), .B1(n_0_0_223), .B2(n_0_59), .C1(n_0_60), 
      .C2(n_0_0_227), .ZN(n_0_0_222));
   OAI21_X1 i_0_0_371 (.A(n_0_0_224), .B1(FIRST_ONE), .B2(Dividend2[4]), 
      .ZN(n_0_0_223));
   NAND2_X1 i_0_0_372 (.A1(n_0_0_316), .A2(FIRST_ONE), .ZN(n_0_0_224));
   OAI21_X1 i_0_0_373 (.A(n_0_0_226), .B1(n_0_0_232), .B2(n_0_0_229), .ZN(
      n_0_0_225));
   AOI22_X1 i_0_0_374 (.A1(n_0_61), .A2(n_0_0_230), .B1(n_0_0_227), .B2(n_0_60), 
      .ZN(n_0_0_226));
   OAI21_X1 i_0_0_375 (.A(n_0_0_228), .B1(FIRST_ONE), .B2(Dividend2[3]), 
      .ZN(n_0_0_227));
   NAND2_X1 i_0_0_376 (.A1(n_0_0_315), .A2(FIRST_ONE), .ZN(n_0_0_228));
   OAI22_X1 i_0_0_377 (.A1(n_0_62), .A2(n_0_0_235), .B1(n_0_0_230), .B2(n_0_61), 
      .ZN(n_0_0_229));
   OAI21_X1 i_0_0_378 (.A(n_0_0_231), .B1(FIRST_ONE), .B2(Dividend2[2]), 
      .ZN(n_0_0_230));
   NAND2_X1 i_0_0_379 (.A1(n_0_0_314), .A2(FIRST_ONE), .ZN(n_0_0_231));
   AOI22_X1 i_0_0_380 (.A1(n_0_62), .A2(n_0_0_235), .B1(n_0_0_233), .B2(n_0_63), 
      .ZN(n_0_0_232));
   OAI21_X1 i_0_0_381 (.A(n_0_0_234), .B1(FIRST_ONE), .B2(Dividend2[0]), 
      .ZN(n_0_0_233));
   NAND2_X1 i_0_0_382 (.A1(n_0_0_312), .A2(FIRST_ONE), .ZN(n_0_0_234));
   OAI21_X1 i_0_0_383 (.A(n_0_0_236), .B1(FIRST_ONE), .B2(Dividend2[1]), 
      .ZN(n_0_0_235));
   NAND2_X1 i_0_0_384 (.A1(n_0_0_313), .A2(FIRST_ONE), .ZN(n_0_0_236));
   NOR2_X1 i_0_0_385 (.A1(n_0_58), .A2(n_0_0_238), .ZN(n_0_0_237));
   OAI21_X1 i_0_0_386 (.A(n_0_0_239), .B1(FIRST_ONE), .B2(Dividend2[5]), 
      .ZN(n_0_0_238));
   NAND2_X1 i_0_0_387 (.A1(n_0_0_317), .A2(FIRST_ONE), .ZN(n_0_0_239));
   AND2_X1 i_0_0_388 (.A1(Index[1]), .A2(Index[0]), .ZN(n_0_0_240));
   NOR4_X1 i_0_0_389 (.A1(n_0_0_283), .A2(n_0_0_241), .A3(n_0_0_279), .A4(rst), 
      .ZN(n_0_216));
   INV_X1 i_0_0_390 (.A(n_0_0_242), .ZN(n_0_0_241));
   OAI21_X1 i_0_0_391 (.A(n_0_0_265), .B1(n_0_0_268), .B2(Divisor[7]), .ZN(
      n_0_0_242));
   NAND2_X1 i_0_0_392 (.A1(n_0_0_276), .A2(n_0_0_243), .ZN(n_0_217));
   AOI21_X1 i_0_0_393 (.A(rst), .B1(n_0_0_244), .B2(n_0_0_328), .ZN(n_0_0_243));
   NOR3_X1 i_0_0_394 (.A1(n_0_0_246), .A2(Index[2]), .A3(Index[3]), .ZN(
      n_0_0_244));
   INV_X1 i_0_0_395 (.A(n_0_0_246), .ZN(n_0_0_245));
   NAND2_X1 i_0_0_396 (.A1(n_0_0_248), .A2(n_0_0_247), .ZN(n_0_0_246));
   NOR2_X1 i_0_0_397 (.A1(Index[1]), .A2(Index[0]), .ZN(n_0_0_247));
   NOR3_X1 i_0_0_398 (.A1(n_0_0_258), .A2(n_0_0_253), .A3(n_0_0_249), .ZN(
      n_0_0_248));
   NAND3_X1 i_0_0_399 (.A1(n_0_0_252), .A2(n_0_0_251), .A3(n_0_0_250), .ZN(
      n_0_0_249));
   NOR2_X1 i_0_0_400 (.A1(Index[21]), .A2(Index[20]), .ZN(n_0_0_250));
   NOR2_X1 i_0_0_401 (.A1(Index[23]), .A2(Index[22]), .ZN(n_0_0_251));
   NOR4_X1 i_0_0_402 (.A1(Index[19]), .A2(Index[18]), .A3(Index[17]), .A4(
      Index[16]), .ZN(n_0_0_252));
   NAND4_X1 i_0_0_403 (.A1(n_0_0_257), .A2(n_0_0_256), .A3(n_0_0_255), .A4(
      n_0_0_254), .ZN(n_0_0_253));
   NOR2_X1 i_0_0_404 (.A1(Index[29]), .A2(Index[28]), .ZN(n_0_0_254));
   NOR2_X1 i_0_0_405 (.A1(Index[31]), .A2(Index[30]), .ZN(n_0_0_255));
   NOR2_X1 i_0_0_406 (.A1(Index[25]), .A2(Index[24]), .ZN(n_0_0_256));
   NOR2_X1 i_0_0_407 (.A1(Index[27]), .A2(Index[26]), .ZN(n_0_0_257));
   NAND3_X1 i_0_0_408 (.A1(n_0_0_261), .A2(n_0_0_260), .A3(n_0_0_259), .ZN(
      n_0_0_258));
   NOR4_X1 i_0_0_409 (.A1(Index[15]), .A2(Index[14]), .A3(Index[13]), .A4(
      Index[12]), .ZN(n_0_0_259));
   NOR4_X1 i_0_0_410 (.A1(Index[11]), .A2(Index[10]), .A3(Index[9]), .A4(
      Index[8]), .ZN(n_0_0_260));
   NOR4_X1 i_0_0_411 (.A1(Index[7]), .A2(Index[6]), .A3(Index[5]), .A4(Index[4]), 
      .ZN(n_0_0_261));
   AOI21_X1 i_0_0_412 (.A(rst), .B1(n_0_0_262), .B2(n_0_2), .ZN(n_0_218));
   NAND3_X1 i_0_0_413 (.A1(n_0_0_264), .A2(n_0_2), .A3(Start), .ZN(n_0_0_262));
   OR2_X1 i_0_0_414 (.A1(n_0_2), .A2(rst), .ZN(n_0_0_263));
   NAND2_X1 i_0_0_415 (.A1(n_0_0_277), .A2(n_0_0_266), .ZN(n_0_0_264));
   NOR2_X1 i_0_0_416 (.A1(n_0_0_266), .A2(n_0_0_276), .ZN(n_0_0_265));
   NOR2_X1 i_0_0_417 (.A1(n_0_0_268), .A2(n_0_0_267), .ZN(n_0_0_266));
   NOR2_X1 i_0_0_418 (.A1(n_0_0_284), .A2(n_0_0_279), .ZN(n_0_0_267));
   NOR2_X1 i_0_0_419 (.A1(n_0_0_305), .A2(n_0_0_269), .ZN(n_0_0_268));
   NAND2_X1 i_0_0_420 (.A1(n_0_0_296), .A2(n_0_0_270), .ZN(n_0_0_269));
   INV_X1 i_0_0_421 (.A(n_0_0_271), .ZN(n_0_0_270));
   NAND3_X1 i_0_0_422 (.A1(n_0_0_293), .A2(n_0_0_338), .A3(n_0_0_339), .ZN(
      n_0_0_271));
   INV_X1 i_0_0_423 (.A(n_0_0_272), .ZN(n_0_219));
   AOI21_X1 i_0_0_424 (.A(rst), .B1(n_0_2), .B2(Start), .ZN(n_0_0_272));
   NOR2_X1 i_0_0_425 (.A1(n_0_0_277), .A2(n_0_0_273), .ZN(n_0_220));
   NAND2_X1 i_0_0_426 (.A1(Start), .A2(n_0_0_275), .ZN(n_0_0_273));
   NOR2_X1 i_0_0_427 (.A1(n_0_0_276), .A2(rst), .ZN(n_0_0_274));
   NOR2_X1 i_0_0_428 (.A1(n_0_0_328), .A2(rst), .ZN(n_0_0_275));
   NAND2_X1 i_0_0_429 (.A1(Start), .A2(n_0_2), .ZN(n_0_0_276));
   OAI211_X1 i_0_0_430 (.A(n_0_0_283), .B(n_0_0_278), .C1(n_0_0_289), .C2(
      n_0_0_305), .ZN(n_0_0_277));
   NOR3_X1 i_0_0_431 (.A1(n_0_0_279), .A2(n_0_0_1), .A3(n_0_0_20), .ZN(n_0_0_278));
   OR3_X1 i_0_0_432 (.A1(n_0_0_281), .A2(n_0_0_280), .A3(Divisor[14]), .ZN(
      n_0_0_279));
   OR2_X1 i_0_0_433 (.A1(Divisor[13]), .A2(Divisor[12]), .ZN(n_0_0_280));
   NAND3_X1 i_0_0_434 (.A1(n_0_0_282), .A2(n_0_0_334), .A3(n_0_0_335), .ZN(
      n_0_0_281));
   NOR2_X1 i_0_0_435 (.A1(Divisor[11]), .A2(Divisor[10]), .ZN(n_0_0_282));
   OR2_X1 i_0_0_436 (.A1(n_0_0_284), .A2(Divisor[7]), .ZN(n_0_0_283));
   OR2_X1 i_0_0_437 (.A1(n_0_0_286), .A2(Divisor[6]), .ZN(n_0_0_284));
   NOR4_X1 i_0_0_438 (.A1(Divisor[7]), .A2(Divisor[6]), .A3(Divisor[5]), 
      .A4(Divisor[4]), .ZN(n_0_0_285));
   OR3_X1 i_0_0_439 (.A1(n_0_0_287), .A2(Divisor[4]), .A3(Divisor[5]), .ZN(
      n_0_0_286));
   NAND3_X1 i_0_0_440 (.A1(n_0_0_288), .A2(n_0_0_329), .A3(n_0_0_330), .ZN(
      n_0_0_287));
   NOR2_X1 i_0_0_441 (.A1(Divisor[3]), .A2(Divisor[2]), .ZN(n_0_0_288));
   AOI211_X1 i_0_0_442 (.A(n_0_0_294), .B(n_0_0_290), .C1(n_0_0_301), .C2(
      n_0_0_298), .ZN(n_0_0_289));
   AOI221_X1 i_0_0_443 (.A(Dividend[14]), .B1(n_0_0_351), .B2(n_0_0_291), 
      .C1(n_0_0_306), .C2(n_0_0_292), .ZN(n_0_0_290));
   AOI21_X1 i_0_0_444 (.A(Dividend[12]), .B1(n_0_0_349), .B2(n_0_0_348), 
      .ZN(n_0_0_291));
   OAI211_X1 i_0_0_445 (.A(n_0_0_345), .B(n_0_0_344), .C1(n_0_0_297), .C2(
      n_0_0_293), .ZN(n_0_0_292));
   NOR2_X1 i_0_0_446 (.A1(Dividend[3]), .A2(Dividend[2]), .ZN(n_0_0_293));
   NOR3_X1 i_0_0_447 (.A1(Dividend[14]), .A2(n_0_0_295), .A3(n_0_0_307), 
      .ZN(n_0_0_294));
   NOR2_X1 i_0_0_448 (.A1(n_0_0_296), .A2(n_0_0_309), .ZN(n_0_0_295));
   NOR3_X1 i_0_0_449 (.A1(n_0_0_297), .A2(Dividend[6]), .A3(Dividend[7]), 
      .ZN(n_0_0_296));
   NAND2_X1 i_0_0_450 (.A1(n_0_0_343), .A2(n_0_0_342), .ZN(n_0_0_297));
   NAND2_X1 i_0_0_451 (.A1(n_0_0_352), .A2(n_0_0_299), .ZN(n_0_0_298));
   OAI21_X1 i_0_0_452 (.A(n_0_0_351), .B1(Dividend[12]), .B2(n_0_0_300), 
      .ZN(n_0_0_299));
   AOI21_X1 i_0_0_453 (.A(Dividend[11]), .B1(n_0_0_348), .B2(Dividend[9]), 
      .ZN(n_0_0_300));
   NAND2_X1 i_0_0_454 (.A1(n_0_0_302), .A2(n_0_0_306), .ZN(n_0_0_301));
   OAI21_X1 i_0_0_455 (.A(n_0_0_345), .B1(Dividend[6]), .B2(n_0_0_303), .ZN(
      n_0_0_302));
   AOI21_X1 i_0_0_456 (.A(Dividend[5]), .B1(n_0_0_342), .B2(n_0_0_304), .ZN(
      n_0_0_303));
   OAI21_X1 i_0_0_457 (.A(n_0_0_341), .B1(n_0_0_339), .B2(Dividend[2]), .ZN(
      n_0_0_304));
   NAND4_X1 i_0_0_458 (.A1(n_0_0_308), .A2(n_0_0_350), .A3(n_0_0_351), .A4(
      n_0_0_352), .ZN(n_0_0_305));
   NOR3_X1 i_0_0_459 (.A1(n_0_0_309), .A2(n_0_0_307), .A3(Dividend[14]), 
      .ZN(n_0_0_306));
   NAND2_X1 i_0_0_460 (.A1(n_0_0_351), .A2(n_0_0_350), .ZN(n_0_0_307));
   INV_X1 i_0_0_461 (.A(n_0_0_309), .ZN(n_0_0_308));
   NAND4_X1 i_0_0_462 (.A1(n_0_0_349), .A2(n_0_0_348), .A3(n_0_0_347), .A4(
      n_0_0_346), .ZN(n_0_0_309));
   INV_X1 i_0_0_463 (.A(n_0_4), .ZN(n_0_0_310));
   INV_X1 i_0_0_464 (.A(n_0_6), .ZN(n_0_0_311));
   INV_X1 i_0_0_465 (.A(addOut[0]), .ZN(n_0_0_312));
   INV_X1 i_0_0_466 (.A(addOut[1]), .ZN(n_0_0_313));
   INV_X1 i_0_0_467 (.A(addOut[2]), .ZN(n_0_0_314));
   INV_X1 i_0_0_468 (.A(addOut[3]), .ZN(n_0_0_315));
   INV_X1 i_0_0_469 (.A(addOut[4]), .ZN(n_0_0_316));
   INV_X1 i_0_0_470 (.A(addOut[5]), .ZN(n_0_0_317));
   INV_X1 i_0_0_471 (.A(addOut[6]), .ZN(n_0_0_318));
   INV_X1 i_0_0_472 (.A(addOut[7]), .ZN(n_0_0_319));
   INV_X1 i_0_0_473 (.A(addOut[8]), .ZN(n_0_0_320));
   INV_X1 i_0_0_474 (.A(addOut[9]), .ZN(n_0_0_321));
   INV_X1 i_0_0_475 (.A(addOut[10]), .ZN(n_0_0_322));
   INV_X1 i_0_0_476 (.A(addOut[11]), .ZN(n_0_0_323));
   INV_X1 i_0_0_477 (.A(addOut[12]), .ZN(n_0_0_324));
   INV_X1 i_0_0_478 (.A(addOut[13]), .ZN(n_0_0_325));
   INV_X1 i_0_0_479 (.A(addOut[14]), .ZN(n_0_0_326));
   INV_X1 i_0_0_480 (.A(addOut[15]), .ZN(n_0_0_327));
   INV_X1 i_0_0_481 (.A(n_0_2), .ZN(n_0_0_328));
   INV_X1 i_0_0_482 (.A(Divisor[0]), .ZN(n_0_0_329));
   INV_X1 i_0_0_483 (.A(Divisor[1]), .ZN(n_0_0_330));
   INV_X1 i_0_0_484 (.A(Divisor[2]), .ZN(n_0_0_331));
   INV_X1 i_0_0_485 (.A(Divisor[5]), .ZN(n_0_0_332));
   INV_X1 i_0_0_486 (.A(Divisor[6]), .ZN(n_0_0_333));
   INV_X1 i_0_0_487 (.A(Divisor[8]), .ZN(n_0_0_334));
   INV_X1 i_0_0_488 (.A(Divisor[9]), .ZN(n_0_0_335));
   INV_X1 i_0_0_489 (.A(Divisor[10]), .ZN(n_0_0_336));
   INV_X1 i_0_0_490 (.A(Divisor[14]), .ZN(n_0_0_337));
   INV_X1 i_0_0_491 (.A(Dividend[0]), .ZN(n_0_0_338));
   INV_X1 i_0_0_492 (.A(Dividend[1]), .ZN(n_0_0_339));
   INV_X1 i_0_0_493 (.A(Dividend[2]), .ZN(n_0_0_340));
   INV_X1 i_0_0_494 (.A(Dividend[3]), .ZN(n_0_0_341));
   INV_X1 i_0_0_495 (.A(Dividend[4]), .ZN(n_0_0_342));
   INV_X1 i_0_0_496 (.A(Dividend[5]), .ZN(n_0_0_343));
   INV_X1 i_0_0_497 (.A(Dividend[6]), .ZN(n_0_0_344));
   INV_X1 i_0_0_498 (.A(Dividend[7]), .ZN(n_0_0_345));
   INV_X1 i_0_0_499 (.A(Dividend[8]), .ZN(n_0_0_346));
   INV_X1 i_0_0_500 (.A(Dividend[9]), .ZN(n_0_0_347));
   INV_X1 i_0_0_501 (.A(Dividend[10]), .ZN(n_0_0_348));
   INV_X1 i_0_0_502 (.A(Dividend[11]), .ZN(n_0_0_349));
   INV_X1 i_0_0_503 (.A(Dividend[12]), .ZN(n_0_0_350));
   INV_X1 i_0_0_504 (.A(Dividend[13]), .ZN(n_0_0_351));
   INV_X1 i_0_0_505 (.A(Dividend[14]), .ZN(n_0_0_352));
   INV_X1 i_0_0_506 (.A(Dividend[15]), .ZN(n_0_0_353));
   INV_X1 i_0_0_507 (.A(Index[0]), .ZN(n_0_0_354));
   INV_X1 i_0_0_508 (.A(Index[3]), .ZN(n_0_0_355));
   INV_X1 i_0_0_509 (.A(n_0_0_263), .ZN(n_0_0_356));
   INV_X1 i_0_0_510 (.A(n_0_0_166), .ZN(n_0_0_357));
   DFF_X1 ERR_reg (.D(n_0_222), .CK(clk), .Q(ERR), .QN());
   DFF_X1 OverFlow_reg (.D(n_0_221), .CK(clk), .Q(OverFlow), .QN());
   MUX2_X1 i_0_1_0 (.A(ERR), .B(n_0_216), .S(n_0_219), .Z(n_0_222));
   MUX2_X1 i_0_1_1 (.A(OverFlow), .B(n_0_220), .S(n_0_219), .Z(n_0_221));
endmodule
