/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 21:06:42 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3318017244 */

module Partial_Full_Adder__0_462(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_458(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_454(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_450(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_446(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_442(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_438(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_434(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_430(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_426(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_422(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_418(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_414(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_410(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_406(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead__0_467(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire c15;
   wire c14;
   wire c13;
   wire c12;
   wire c11;
   wire c10;
   wire c9;
   wire c8;
   wire c7;
   wire c6;
   wire c5;
   wire c4;
   wire c3;
   wire c2;

   Partial_Full_Adder__0_462 PFA2 (.A(A[1]), .B(), .Cin(A[0]), .S(S[1]), .P(), 
      .G());
   Partial_Full_Adder__0_458 PFA3 (.A(A[2]), .B(), .Cin(c2), .S(S[2]), .P(), 
      .G());
   Partial_Full_Adder__0_454 PFA4 (.A(A[3]), .B(), .Cin(c3), .S(S[3]), .P(), 
      .G());
   Partial_Full_Adder__0_450 PFA5 (.A(A[4]), .B(), .Cin(c4), .S(S[4]), .P(), 
      .G());
   Partial_Full_Adder__0_446 PFA6 (.A(A[5]), .B(), .Cin(c5), .S(S[5]), .P(), 
      .G());
   Partial_Full_Adder__0_442 PFA7 (.A(A[6]), .B(), .Cin(c6), .S(S[6]), .P(), 
      .G());
   Partial_Full_Adder__0_438 PFA8 (.A(A[7]), .B(), .Cin(c7), .S(S[7]), .P(), 
      .G());
   Partial_Full_Adder__0_434 PFA9 (.A(A[8]), .B(), .Cin(c8), .S(S[8]), .P(), 
      .G());
   Partial_Full_Adder__0_430 PFA10 (.A(A[9]), .B(), .Cin(c9), .S(S[9]), .P(), 
      .G());
   Partial_Full_Adder__0_426 PFA11 (.A(A[10]), .B(), .Cin(c10), .S(S[10]), .P(), 
      .G());
   Partial_Full_Adder__0_422 PFA12 (.A(A[11]), .B(), .Cin(c11), .S(S[11]), .P(), 
      .G());
   Partial_Full_Adder__0_418 PFA13 (.A(A[12]), .B(), .Cin(c12), .S(S[12]), .P(), 
      .G());
   Partial_Full_Adder__0_414 PFA14 (.A(A[13]), .B(), .Cin(c13), .S(S[13]), .P(), 
      .G());
   Partial_Full_Adder__0_410 PFA15 (.A(A[14]), .B(), .Cin(c14), .S(S[14]), .P(), 
      .G());
   Partial_Full_Adder__0_406 PFA16 (.A(A[15]), .B(), .Cin(c15), .S(S[15]), .P(), 
      .G());
   AND2_X1 i_0_0 (.A1(A[14]), .A2(c14), .ZN(c15));
   AND2_X1 i_0_1 (.A1(A[13]), .A2(c13), .ZN(c14));
   AND2_X1 i_0_2 (.A1(A[12]), .A2(c12), .ZN(c13));
   AND2_X1 i_0_3 (.A1(A[11]), .A2(c11), .ZN(c12));
   AND2_X1 i_0_4 (.A1(A[10]), .A2(c10), .ZN(c11));
   AND2_X1 i_0_5 (.A1(A[9]), .A2(c9), .ZN(c10));
   AND2_X1 i_0_6 (.A1(A[8]), .A2(c8), .ZN(c9));
   AND2_X1 i_0_7 (.A1(A[7]), .A2(c7), .ZN(c8));
   AND2_X1 i_0_8 (.A1(A[6]), .A2(c6), .ZN(c7));
   AND2_X1 i_0_9 (.A1(A[5]), .A2(c5), .ZN(c6));
   AND2_X1 i_0_10 (.A1(A[4]), .A2(c4), .ZN(c5));
   AND2_X1 i_0_11 (.A1(A[3]), .A2(c3), .ZN(c4));
   AND2_X1 i_0_12 (.A1(A[2]), .A2(c2), .ZN(c3));
   AND2_X1 i_0_13 (.A1(A[0]), .A2(A[1]), .ZN(c2));
endmodule

module Partial_Full_Adder__0_547(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_543(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_539(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_535(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_531(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_527(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_523(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_519(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_515(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_511(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_507(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_503(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_499(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_495(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_491(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_487(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead__0_548(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire c1;
   wire c15;
   wire n_0_0;
   wire c14;
   wire n_0_1;
   wire c13;
   wire n_0_2;
   wire c12;
   wire n_0_3;
   wire c11;
   wire n_0_4;
   wire c10;
   wire n_0_5;
   wire c9;
   wire n_0_6;
   wire c8;
   wire n_0_7;
   wire c7;
   wire n_0_8;
   wire c6;
   wire n_0_9;
   wire c5;
   wire n_0_10;
   wire c4;
   wire n_0_11;
   wire c3;
   wire n_0_12;
   wire c2;
   wire n_0_13;

   Partial_Full_Adder__0_547 PFA1 (.A(A[0]), .B(B[0]), .Cin(), .S(S[0]), .P(), 
      .G(c1));
   Partial_Full_Adder__0_543 PFA2 (.A(A[1]), .B(B[1]), .Cin(c1), .S(S[1]), 
      .P(n_1), .G(n_0));
   Partial_Full_Adder__0_539 PFA3 (.A(A[2]), .B(B[2]), .Cin(c2), .S(S[2]), 
      .P(n_3), .G(n_2));
   Partial_Full_Adder__0_535 PFA4 (.A(A[3]), .B(B[3]), .Cin(c3), .S(S[3]), 
      .P(n_5), .G(n_4));
   Partial_Full_Adder__0_531 PFA5 (.A(A[4]), .B(B[4]), .Cin(c4), .S(S[4]), 
      .P(n_7), .G(n_6));
   Partial_Full_Adder__0_527 PFA6 (.A(A[5]), .B(B[5]), .Cin(c5), .S(S[5]), 
      .P(n_9), .G(n_8));
   Partial_Full_Adder__0_523 PFA7 (.A(A[6]), .B(B[6]), .Cin(c6), .S(S[6]), 
      .P(n_11), .G(n_10));
   Partial_Full_Adder__0_519 PFA8 (.A(A[7]), .B(B[7]), .Cin(c7), .S(S[7]), 
      .P(n_13), .G(n_12));
   Partial_Full_Adder__0_515 PFA9 (.A(A[8]), .B(B[8]), .Cin(c8), .S(S[8]), 
      .P(n_15), .G(n_14));
   Partial_Full_Adder__0_511 PFA10 (.A(A[9]), .B(B[9]), .Cin(c9), .S(S[9]), 
      .P(n_17), .G(n_16));
   Partial_Full_Adder__0_507 PFA11 (.A(A[10]), .B(B[10]), .Cin(c10), .S(S[10]), 
      .P(n_19), .G(n_18));
   Partial_Full_Adder__0_503 PFA12 (.A(A[11]), .B(B[11]), .Cin(c11), .S(S[11]), 
      .P(n_21), .G(n_20));
   Partial_Full_Adder__0_499 PFA13 (.A(A[12]), .B(B[12]), .Cin(c12), .S(S[12]), 
      .P(n_23), .G(n_22));
   Partial_Full_Adder__0_495 PFA14 (.A(A[13]), .B(B[13]), .Cin(c13), .S(S[13]), 
      .P(n_25), .G(n_24));
   Partial_Full_Adder__0_491 PFA15 (.A(A[14]), .B(B[14]), .Cin(c14), .S(S[14]), 
      .P(n_27), .G(n_26));
   Partial_Full_Adder__0_487 PFA16 (.A(A[15]), .B(B[15]), .Cin(c15), .S(S[15]), 
      .P(), .G());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(c15));
   AOI21_X1 i_0_1 (.A(n_26), .B1(n_27), .B2(c14), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(c14));
   AOI21_X1 i_0_3 (.A(n_24), .B1(n_25), .B2(c13), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(c13));
   AOI21_X1 i_0_5 (.A(n_22), .B1(n_23), .B2(c12), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(c12));
   AOI21_X1 i_0_7 (.A(n_20), .B1(n_21), .B2(c11), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(c11));
   AOI21_X1 i_0_9 (.A(n_18), .B1(n_19), .B2(c10), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(c10));
   AOI21_X1 i_0_11 (.A(n_16), .B1(n_17), .B2(c9), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(c9));
   AOI21_X1 i_0_13 (.A(n_14), .B1(n_15), .B2(c8), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(c8));
   AOI21_X1 i_0_15 (.A(n_12), .B1(n_13), .B2(c7), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(c7));
   AOI21_X1 i_0_17 (.A(n_10), .B1(n_11), .B2(c6), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(c6));
   AOI21_X1 i_0_19 (.A(n_8), .B1(n_9), .B2(c5), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(c5));
   AOI21_X1 i_0_21 (.A(n_6), .B1(n_7), .B2(c4), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(c4));
   AOI21_X1 i_0_23 (.A(n_4), .B1(n_5), .B2(c3), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(c3));
   AOI21_X1 i_0_25 (.A(n_2), .B1(n_3), .B2(c2), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(c2));
   AOI21_X1 i_0_27 (.A(n_0), .B1(c1), .B2(n_1), .ZN(n_0_13));
endmodule

module Partial_Full_Adder__0_628(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_624(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_620(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_616(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_612(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_608(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_604(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_600(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_596(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_592(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_588(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_584(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_580(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_576(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_572(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_568(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead__0_629(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire c1;
   wire c15;
   wire n_0_0;
   wire c14;
   wire n_0_1;
   wire c13;
   wire n_0_2;
   wire c12;
   wire n_0_3;
   wire c11;
   wire n_0_4;
   wire c10;
   wire n_0_5;
   wire c9;
   wire n_0_6;
   wire c8;
   wire n_0_7;
   wire c7;
   wire n_0_8;
   wire c6;
   wire n_0_9;
   wire c5;
   wire n_0_10;
   wire c4;
   wire n_0_11;
   wire c3;
   wire n_0_12;
   wire c2;
   wire n_0_13;

   Partial_Full_Adder__0_628 PFA1 (.A(A[0]), .B(B[0]), .Cin(), .S(S[0]), .P(), 
      .G(c1));
   Partial_Full_Adder__0_624 PFA2 (.A(A[1]), .B(B[1]), .Cin(c1), .S(S[1]), 
      .P(n_1), .G(n_0));
   Partial_Full_Adder__0_620 PFA3 (.A(A[2]), .B(B[2]), .Cin(c2), .S(S[2]), 
      .P(n_3), .G(n_2));
   Partial_Full_Adder__0_616 PFA4 (.A(A[3]), .B(B[3]), .Cin(c3), .S(S[3]), 
      .P(n_5), .G(n_4));
   Partial_Full_Adder__0_612 PFA5 (.A(A[4]), .B(B[4]), .Cin(c4), .S(S[4]), 
      .P(n_7), .G(n_6));
   Partial_Full_Adder__0_608 PFA6 (.A(A[5]), .B(B[5]), .Cin(c5), .S(S[5]), 
      .P(n_9), .G(n_8));
   Partial_Full_Adder__0_604 PFA7 (.A(A[6]), .B(B[6]), .Cin(c6), .S(S[6]), 
      .P(n_11), .G(n_10));
   Partial_Full_Adder__0_600 PFA8 (.A(A[7]), .B(B[7]), .Cin(c7), .S(S[7]), 
      .P(n_13), .G(n_12));
   Partial_Full_Adder__0_596 PFA9 (.A(A[8]), .B(B[8]), .Cin(c8), .S(S[8]), 
      .P(n_15), .G(n_14));
   Partial_Full_Adder__0_592 PFA10 (.A(A[9]), .B(B[9]), .Cin(c9), .S(S[9]), 
      .P(n_17), .G(n_16));
   Partial_Full_Adder__0_588 PFA11 (.A(A[10]), .B(B[10]), .Cin(c10), .S(S[10]), 
      .P(n_19), .G(n_18));
   Partial_Full_Adder__0_584 PFA12 (.A(A[11]), .B(B[11]), .Cin(c11), .S(S[11]), 
      .P(n_21), .G(n_20));
   Partial_Full_Adder__0_580 PFA13 (.A(A[12]), .B(B[12]), .Cin(c12), .S(S[12]), 
      .P(n_23), .G(n_22));
   Partial_Full_Adder__0_576 PFA14 (.A(A[13]), .B(B[13]), .Cin(c13), .S(S[13]), 
      .P(n_25), .G(n_24));
   Partial_Full_Adder__0_572 PFA15 (.A(A[14]), .B(B[14]), .Cin(c14), .S(S[14]), 
      .P(n_27), .G(n_26));
   Partial_Full_Adder__0_568 PFA16 (.A(A[15]), .B(B[15]), .Cin(c15), .S(S[15]), 
      .P(), .G());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(c15));
   AOI21_X1 i_0_1 (.A(n_26), .B1(n_27), .B2(c14), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(c14));
   AOI21_X1 i_0_3 (.A(n_24), .B1(n_25), .B2(c13), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(c13));
   AOI21_X1 i_0_5 (.A(n_22), .B1(n_23), .B2(c12), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(c12));
   AOI21_X1 i_0_7 (.A(n_20), .B1(n_21), .B2(c11), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(c11));
   AOI21_X1 i_0_9 (.A(n_18), .B1(n_19), .B2(c10), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(c10));
   AOI21_X1 i_0_11 (.A(n_16), .B1(n_17), .B2(c9), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(c9));
   AOI21_X1 i_0_13 (.A(n_14), .B1(n_15), .B2(c8), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(c8));
   AOI21_X1 i_0_15 (.A(n_12), .B1(n_13), .B2(c7), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(c7));
   AOI21_X1 i_0_17 (.A(n_10), .B1(n_11), .B2(c6), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(c6));
   AOI21_X1 i_0_19 (.A(n_8), .B1(n_9), .B2(c5), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(c5));
   AOI21_X1 i_0_21 (.A(n_6), .B1(n_7), .B2(c4), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(c4));
   AOI21_X1 i_0_23 (.A(n_4), .B1(n_5), .B2(c3), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(c3));
   AOI21_X1 i_0_25 (.A(n_2), .B1(n_3), .B2(c2), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(c2));
   AOI21_X1 i_0_27 (.A(n_0), .B1(c1), .B2(n_1), .ZN(n_0_13));
endmodule

module flipflop__0_835(D, load, Clk, Q, rst);
   input D;
   input load;
   input Clk;
   output Q;
   input rst;

   DFFR_X1 Q_reg (.D(n_0), .RN(D), .CK(n_1), .Q(Q), .QN());
   MUX2_X1 Q_reg_enable_mux_0 (.A(Q), .B(D), .S(load), .Z(n_0));
   INV_X1 i_0_0 (.A(Clk), .ZN(n_1));
endmodule

module flipflop(D, load, Clk, Q, rst);
   input D;
   input load;
   input Clk;
   output Q;
   input rst;

   DFFR_X1 Q_reg (.D(n_0), .RN(n_2), .CK(n_1), .Q(Q), .QN());
   MUX2_X1 Q_reg_enable_mux_0 (.A(Q), .B(D), .S(load), .Z(n_0));
   INV_X1 i_0_0 (.A(Clk), .ZN(n_1));
   INV_X1 i_1_0 (.A(rst), .ZN(n_2));
endmodule

module Partial_Full_Adder__0_385(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   INV_X1 i_3 (.A(P), .ZN(S));
   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_381(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_377(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_373(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_369(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_365(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_361(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_357(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_353(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_349(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_345(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_341(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_337(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_333(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_329(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_325(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead__0_386(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire G;
   wire P;
   wire c15;
   wire n_0_0;
   wire c14;
   wire n_0_1;
   wire c13;
   wire n_0_2;
   wire c12;
   wire n_0_3;
   wire c11;
   wire n_0_4;
   wire c10;
   wire n_0_5;
   wire c9;
   wire n_0_6;
   wire c8;
   wire n_0_7;
   wire c7;
   wire n_0_8;
   wire c6;
   wire n_0_9;
   wire c5;
   wire n_0_10;
   wire c4;
   wire n_0_11;
   wire c3;
   wire n_0_12;
   wire c2;
   wire n_0_13;
   wire c1;

   Partial_Full_Adder__0_385 PFA1 (.A(A[0]), .B(B[0]), .Cin(), .S(S[0]), 
      .P(P), .G(G));
   Partial_Full_Adder__0_381 PFA2 (.A(A[1]), .B(B[1]), .Cin(c1), .S(S[1]), 
      .P(n_1), .G(n_0));
   Partial_Full_Adder__0_377 PFA3 (.A(A[2]), .B(B[2]), .Cin(c2), .S(S[2]), 
      .P(n_3), .G(n_2));
   Partial_Full_Adder__0_373 PFA4 (.A(A[3]), .B(B[3]), .Cin(c3), .S(S[3]), 
      .P(n_5), .G(n_4));
   Partial_Full_Adder__0_369 PFA5 (.A(A[4]), .B(B[4]), .Cin(c4), .S(S[4]), 
      .P(n_7), .G(n_6));
   Partial_Full_Adder__0_365 PFA6 (.A(A[5]), .B(B[5]), .Cin(c5), .S(S[5]), 
      .P(n_9), .G(n_8));
   Partial_Full_Adder__0_361 PFA7 (.A(A[6]), .B(B[6]), .Cin(c6), .S(S[6]), 
      .P(n_11), .G(n_10));
   Partial_Full_Adder__0_357 PFA8 (.A(A[7]), .B(B[7]), .Cin(c7), .S(S[7]), 
      .P(n_13), .G(n_12));
   Partial_Full_Adder__0_353 PFA9 (.A(A[8]), .B(B[8]), .Cin(c8), .S(S[8]), 
      .P(n_15), .G(n_14));
   Partial_Full_Adder__0_349 PFA10 (.A(A[9]), .B(B[9]), .Cin(c9), .S(S[9]), 
      .P(n_17), .G(n_16));
   Partial_Full_Adder__0_345 PFA11 (.A(A[10]), .B(B[10]), .Cin(c10), .S(S[10]), 
      .P(n_19), .G(n_18));
   Partial_Full_Adder__0_341 PFA12 (.A(A[11]), .B(B[11]), .Cin(c11), .S(S[11]), 
      .P(n_21), .G(n_20));
   Partial_Full_Adder__0_337 PFA13 (.A(A[12]), .B(B[12]), .Cin(c12), .S(S[12]), 
      .P(n_23), .G(n_22));
   Partial_Full_Adder__0_333 PFA14 (.A(A[13]), .B(B[13]), .Cin(c13), .S(S[13]), 
      .P(n_25), .G(n_24));
   Partial_Full_Adder__0_329 PFA15 (.A(A[14]), .B(B[14]), .Cin(c14), .S(S[14]), 
      .P(n_27), .G(n_26));
   Partial_Full_Adder__0_325 PFA16 (.A(A[15]), .B(B[15]), .Cin(c15), .S(S[15]), 
      .P(), .G());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(c15));
   AOI21_X1 i_0_1 (.A(n_26), .B1(n_27), .B2(c14), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(c14));
   AOI21_X1 i_0_3 (.A(n_24), .B1(n_25), .B2(c13), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(c13));
   AOI21_X1 i_0_5 (.A(n_22), .B1(n_23), .B2(c12), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(c12));
   AOI21_X1 i_0_7 (.A(n_20), .B1(n_21), .B2(c11), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(c11));
   AOI21_X1 i_0_9 (.A(n_18), .B1(n_19), .B2(c10), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(c10));
   AOI21_X1 i_0_11 (.A(n_16), .B1(n_17), .B2(c9), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(c9));
   AOI21_X1 i_0_13 (.A(n_14), .B1(n_15), .B2(c8), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(c8));
   AOI21_X1 i_0_15 (.A(n_12), .B1(n_13), .B2(c7), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(c7));
   AOI21_X1 i_0_17 (.A(n_10), .B1(n_11), .B2(c6), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(c6));
   AOI21_X1 i_0_19 (.A(n_8), .B1(n_9), .B2(c5), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(c5));
   AOI21_X1 i_0_21 (.A(n_6), .B1(n_7), .B2(c4), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(c4));
   AOI21_X1 i_0_23 (.A(n_4), .B1(n_5), .B2(c3), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(c3));
   AOI21_X1 i_0_25 (.A(n_2), .B1(n_3), .B2(c2), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(c2));
   AOI21_X1 i_0_27 (.A(n_0), .B1(n_1), .B2(c1), .ZN(n_0_13));
   OR2_X1 i_0_28 (.A1(P), .A2(G), .ZN(c1));
endmodule

module datapath__0_59(Index, p_0);
   input [31:0]Index;
   output [31:0]p_0;

   INV_X1 i_0 (.A(Index[0]), .ZN(p_0[0]));
   XNOR2_X1 i_1 (.A(Index[1]), .B(Index[0]), .ZN(p_0[1]));
   OR2_X1 i_2 (.A1(Index[1]), .A2(Index[0]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(Index[2]), .B(n_0), .ZN(p_0[2]));
   OR2_X1 i_4 (.A1(Index[2]), .A2(n_0), .ZN(n_1));
   XNOR2_X1 i_5 (.A(Index[3]), .B(n_1), .ZN(p_0[3]));
   OR2_X1 i_6 (.A1(Index[3]), .A2(n_1), .ZN(n_2));
   XNOR2_X1 i_7 (.A(Index[4]), .B(n_2), .ZN(p_0[4]));
   OR2_X1 i_8 (.A1(Index[4]), .A2(n_2), .ZN(n_3));
   XNOR2_X1 i_9 (.A(Index[5]), .B(n_3), .ZN(p_0[5]));
   OR2_X1 i_10 (.A1(Index[5]), .A2(n_3), .ZN(n_4));
   XNOR2_X1 i_11 (.A(Index[6]), .B(n_4), .ZN(p_0[6]));
   OR2_X1 i_12 (.A1(Index[6]), .A2(n_4), .ZN(n_5));
   XNOR2_X1 i_13 (.A(Index[7]), .B(n_5), .ZN(p_0[7]));
   OR2_X1 i_14 (.A1(Index[7]), .A2(n_5), .ZN(n_6));
   XNOR2_X1 i_15 (.A(Index[8]), .B(n_6), .ZN(p_0[8]));
   OR2_X1 i_16 (.A1(Index[8]), .A2(n_6), .ZN(n_7));
   XNOR2_X1 i_17 (.A(Index[9]), .B(n_7), .ZN(p_0[9]));
   OR2_X1 i_18 (.A1(Index[9]), .A2(n_7), .ZN(n_8));
   XNOR2_X1 i_19 (.A(Index[10]), .B(n_8), .ZN(p_0[10]));
   OR2_X1 i_20 (.A1(Index[10]), .A2(n_8), .ZN(n_9));
   XNOR2_X1 i_21 (.A(Index[11]), .B(n_9), .ZN(p_0[11]));
   OR2_X1 i_22 (.A1(Index[11]), .A2(n_9), .ZN(n_10));
   XNOR2_X1 i_23 (.A(Index[12]), .B(n_10), .ZN(p_0[12]));
   OR2_X1 i_24 (.A1(Index[12]), .A2(n_10), .ZN(n_11));
   XNOR2_X1 i_25 (.A(Index[13]), .B(n_11), .ZN(p_0[13]));
   OR2_X1 i_26 (.A1(Index[13]), .A2(n_11), .ZN(n_12));
   XNOR2_X1 i_27 (.A(Index[14]), .B(n_12), .ZN(p_0[14]));
   OR2_X1 i_28 (.A1(Index[14]), .A2(n_12), .ZN(n_13));
   XNOR2_X1 i_29 (.A(Index[15]), .B(n_13), .ZN(p_0[15]));
   OR2_X1 i_30 (.A1(Index[15]), .A2(n_13), .ZN(n_14));
   XNOR2_X1 i_31 (.A(Index[16]), .B(n_14), .ZN(p_0[16]));
   OR2_X1 i_32 (.A1(Index[16]), .A2(n_14), .ZN(n_15));
   XNOR2_X1 i_33 (.A(Index[17]), .B(n_15), .ZN(p_0[17]));
   OR2_X1 i_34 (.A1(Index[17]), .A2(n_15), .ZN(n_16));
   XNOR2_X1 i_35 (.A(Index[18]), .B(n_16), .ZN(p_0[18]));
   OR2_X1 i_36 (.A1(Index[18]), .A2(n_16), .ZN(n_17));
   XNOR2_X1 i_37 (.A(Index[19]), .B(n_17), .ZN(p_0[19]));
   OR2_X1 i_38 (.A1(Index[19]), .A2(n_17), .ZN(n_18));
   XNOR2_X1 i_39 (.A(Index[20]), .B(n_18), .ZN(p_0[20]));
   OR2_X1 i_40 (.A1(Index[20]), .A2(n_18), .ZN(n_19));
   XNOR2_X1 i_41 (.A(Index[21]), .B(n_19), .ZN(p_0[21]));
   OR2_X1 i_42 (.A1(Index[21]), .A2(n_19), .ZN(n_20));
   XNOR2_X1 i_43 (.A(Index[22]), .B(n_20), .ZN(p_0[22]));
   OR2_X1 i_44 (.A1(Index[22]), .A2(n_20), .ZN(n_21));
   XNOR2_X1 i_45 (.A(Index[23]), .B(n_21), .ZN(p_0[23]));
   OR2_X1 i_46 (.A1(Index[23]), .A2(n_21), .ZN(n_22));
   XNOR2_X1 i_47 (.A(Index[24]), .B(n_22), .ZN(p_0[24]));
   OR2_X1 i_48 (.A1(Index[24]), .A2(n_22), .ZN(n_23));
   XNOR2_X1 i_49 (.A(Index[25]), .B(n_23), .ZN(p_0[25]));
   OR2_X1 i_50 (.A1(Index[25]), .A2(n_23), .ZN(n_24));
   XNOR2_X1 i_51 (.A(Index[26]), .B(n_24), .ZN(p_0[26]));
   OR2_X1 i_52 (.A1(Index[26]), .A2(n_24), .ZN(n_25));
   XNOR2_X1 i_53 (.A(Index[27]), .B(n_25), .ZN(p_0[27]));
   OR2_X1 i_54 (.A1(Index[27]), .A2(n_25), .ZN(n_26));
   XNOR2_X1 i_55 (.A(Index[28]), .B(n_26), .ZN(p_0[28]));
   OR2_X1 i_56 (.A1(Index[28]), .A2(n_26), .ZN(n_27));
   XNOR2_X1 i_57 (.A(Index[29]), .B(n_27), .ZN(p_0[29]));
   OR2_X1 i_58 (.A1(Index[29]), .A2(n_27), .ZN(n_28));
   XNOR2_X1 i_59 (.A(Index[30]), .B(n_28), .ZN(p_0[30]));
   OR2_X1 i_60 (.A1(Index[30]), .A2(n_28), .ZN(n_29));
   XNOR2_X1 i_61 (.A(Index[31]), .B(n_29), .ZN(p_0[31]));
endmodule

module fixed_division(Dividend, Divisor, Reset, clk, Start, Quotient, ERR, Done, 
      OverFlow);
   input [15:0]Dividend;
   input [15:0]Divisor;
   input Reset;
   input clk;
   input Start;
   output [15:0]Quotient;
   output ERR;
   output Done;
   output OverFlow;

   wire [15:0]addOut;
   wire [15:0]add2;
   wire [15:0]add1;
   wire n_0_19__0;
   wire n_0_20;
   wire n_0_0;
   wire n_0_1;
   wire n_0_16;
   wire n_0_2;
   wire n_0_14__0;
   wire n_0_3;
   wire n_0_15;
   wire n_0_4__0;
   wire n_0_13;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9__0;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_17;
   wire n_0_18;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24__0;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29__0;
   wire n_0_30;
   wire n_0_31;
   wire [15:0]Dividend2;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34__0;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39__0;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44__0;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49__0;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54__0;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59__0;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64__0;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69__0;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74__0;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire [15:0]QuotientVar;
   wire [31:0]Index;
   wire n_0_123;
   wire FIRST_ONE;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_4__1;
   wire n_0_9__1;
   wire n_0_14__1;
   wire n_0_19__1;
   wire n_0_24__1;
   wire n_0_29__1;
   wire n_0_34__1;
   wire n_0_39__1;
   wire n_0_44__1;
   wire n_0_49__1;
   wire n_0_54__1;
   wire n_0_59__1;
   wire n_0_64__1;
   wire n_0_69__1;
   wire n_0_74__1;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;

   Carry_Look_Ahead__0_386 u1 (.A(add1), .B(add2), .Cin(), .S(addOut));
   DLH_X1 Done_reg (.D(n_196), .G(n_194), .Q(Done));
   DLH_X1 \Quotient_reg[15]  (.D(n_193), .G(n_177), .Q(Quotient[15]));
   DLH_X1 \Quotient_reg[14]  (.D(n_192), .G(n_177), .Q(Quotient[14]));
   DLH_X1 \Quotient_reg[13]  (.D(n_191), .G(n_177), .Q(Quotient[13]));
   DLH_X1 \Quotient_reg[12]  (.D(n_190), .G(n_177), .Q(Quotient[12]));
   DLH_X1 \Quotient_reg[11]  (.D(n_189), .G(n_177), .Q(Quotient[11]));
   DLH_X1 \Quotient_reg[10]  (.D(n_188), .G(n_177), .Q(Quotient[10]));
   DLH_X1 \Quotient_reg[9]  (.D(n_187), .G(n_177), .Q(Quotient[9]));
   DLH_X1 \Quotient_reg[8]  (.D(n_186), .G(n_177), .Q(Quotient[8]));
   DLH_X1 \Quotient_reg[7]  (.D(n_185), .G(n_177), .Q(Quotient[7]));
   DLH_X1 \Quotient_reg[6]  (.D(n_184), .G(n_177), .Q(Quotient[6]));
   DLH_X1 \Quotient_reg[5]  (.D(n_183), .G(n_177), .Q(Quotient[5]));
   DLH_X1 \Quotient_reg[4]  (.D(n_182), .G(n_177), .Q(Quotient[4]));
   DLH_X1 \Quotient_reg[3]  (.D(n_181), .G(n_177), .Q(Quotient[3]));
   DLH_X1 \Quotient_reg[2]  (.D(n_180), .G(n_177), .Q(Quotient[2]));
   DLH_X1 \Quotient_reg[1]  (.D(n_179), .G(n_177), .Q(Quotient[1]));
   DLH_X1 \Quotient_reg[0]  (.D(n_178), .G(n_177), .Q(Quotient[0]));
   DLH_X1 \add2_reg[15]  (.D(n_0_74__1), .G(n_176), .Q(add2[15]));
   DLH_X1 \add2_reg[14]  (.D(n_0_69__1), .G(n_176), .Q(add2[14]));
   DLH_X1 \add2_reg[13]  (.D(n_0_64__1), .G(n_176), .Q(add2[13]));
   DLH_X1 \add2_reg[12]  (.D(n_0_59__1), .G(n_176), .Q(add2[12]));
   DLH_X1 \add2_reg[11]  (.D(n_0_54__1), .G(n_176), .Q(add2[11]));
   DLH_X1 \add2_reg[10]  (.D(n_0_49__1), .G(n_176), .Q(add2[10]));
   DLH_X1 \add2_reg[9]  (.D(n_0_44__1), .G(n_176), .Q(add2[9]));
   DLH_X1 \add2_reg[8]  (.D(n_0_39__1), .G(n_176), .Q(add2[8]));
   DLH_X1 \add2_reg[7]  (.D(n_0_34__1), .G(n_176), .Q(add2[7]));
   DLH_X1 \add2_reg[6]  (.D(n_0_29__1), .G(n_176), .Q(add2[6]));
   DLH_X1 \add2_reg[5]  (.D(n_0_24__1), .G(n_176), .Q(add2[5]));
   DLH_X1 \add2_reg[4]  (.D(n_0_19__1), .G(n_176), .Q(add2[4]));
   DLH_X1 \add2_reg[3]  (.D(n_0_14__1), .G(n_176), .Q(add2[3]));
   DLH_X1 \add2_reg[2]  (.D(n_0_9__1), .G(n_176), .Q(add2[2]));
   DLH_X1 \add2_reg[1]  (.D(n_0_4__1), .G(n_176), .Q(add2[1]));
   DLH_X1 \add2_reg[0]  (.D(n_213), .G(n_176), .Q(add2[0]));
   DLH_X1 \add1_reg[15]  (.D(n_212), .G(n_176), .Q(add1[15]));
   DLH_X1 \add1_reg[14]  (.D(n_211), .G(n_176), .Q(add1[14]));
   DLH_X1 \add1_reg[13]  (.D(n_210), .G(n_176), .Q(add1[13]));
   DLH_X1 \add1_reg[12]  (.D(n_209), .G(n_176), .Q(add1[12]));
   DLH_X1 \add1_reg[11]  (.D(n_208), .G(n_176), .Q(add1[11]));
   DLH_X1 \add1_reg[10]  (.D(n_207), .G(n_176), .Q(add1[10]));
   DLH_X1 \add1_reg[9]  (.D(n_206), .G(n_176), .Q(add1[9]));
   DLH_X1 \add1_reg[8]  (.D(n_205), .G(n_176), .Q(add1[8]));
   DLH_X1 \add1_reg[7]  (.D(n_204), .G(n_176), .Q(add1[7]));
   DLH_X1 \add1_reg[6]  (.D(n_203), .G(n_176), .Q(add1[6]));
   DLH_X1 \add1_reg[5]  (.D(n_202), .G(n_176), .Q(add1[5]));
   DLH_X1 \add1_reg[4]  (.D(n_201), .G(n_176), .Q(add1[4]));
   DLH_X1 \add1_reg[3]  (.D(n_200), .G(n_176), .Q(add1[3]));
   DLH_X1 \add1_reg[2]  (.D(n_199), .G(n_176), .Q(add1[2]));
   DLH_X1 \add1_reg[1]  (.D(n_198), .G(n_176), .Q(add1[1]));
   DLH_X1 \add1_reg[0]  (.D(n_197), .G(n_176), .Q(add1[0]));
   DLH_X1 Done_bit_reg (.D(n_175), .G(n_174), .Q(n_0));
   DLH_X1 \Index_reg[31]  (.D(Index[31]), .G(n_195), .Q(n_1));
   DLH_X1 \Index_reg[30]  (.D(Index[30]), .G(n_195), .Q(n_2));
   DLH_X1 \Index_reg[29]  (.D(Index[29]), .G(n_195), .Q(n_3));
   DLH_X1 \Index_reg[28]  (.D(Index[28]), .G(n_195), .Q(n_4));
   DLH_X1 \Index_reg[27]  (.D(Index[27]), .G(n_195), .Q(n_5));
   DLH_X1 \Index_reg[26]  (.D(Index[26]), .G(n_195), .Q(n_6));
   DLH_X1 \Index_reg[25]  (.D(Index[25]), .G(n_195), .Q(n_7));
   DLH_X1 \Index_reg[24]  (.D(Index[24]), .G(n_195), .Q(n_8));
   DLH_X1 \Index_reg[23]  (.D(Index[23]), .G(n_195), .Q(n_9));
   DLH_X1 \Index_reg[22]  (.D(Index[22]), .G(n_195), .Q(n_10));
   DLH_X1 \Index_reg[21]  (.D(Index[21]), .G(n_195), .Q(n_11));
   DLH_X1 \Index_reg[20]  (.D(Index[20]), .G(n_195), .Q(n_12));
   DLH_X1 \Index_reg[19]  (.D(Index[19]), .G(n_195), .Q(n_13));
   DLH_X1 \Index_reg[18]  (.D(Index[18]), .G(n_195), .Q(n_14));
   DLH_X1 \Index_reg[17]  (.D(Index[17]), .G(n_195), .Q(n_15));
   DLH_X1 \Index_reg[16]  (.D(Index[16]), .G(n_195), .Q(n_16));
   DLH_X1 \Index_reg[15]  (.D(Index[15]), .G(n_195), .Q(n_17));
   DLH_X1 \Index_reg[14]  (.D(Index[14]), .G(n_195), .Q(n_18));
   DLH_X1 \Index_reg[13]  (.D(Index[13]), .G(n_195), .Q(n_19));
   DLH_X1 \Index_reg[12]  (.D(Index[12]), .G(n_195), .Q(n_20));
   DLH_X1 \Index_reg[11]  (.D(Index[11]), .G(n_195), .Q(n_21));
   DLH_X1 \Index_reg[10]  (.D(Index[10]), .G(n_195), .Q(n_22));
   DLH_X1 \Index_reg[9]  (.D(Index[9]), .G(n_195), .Q(n_23));
   DLH_X1 \Index_reg[8]  (.D(Index[8]), .G(n_195), .Q(n_24));
   DLH_X1 \Index_reg[7]  (.D(Index[7]), .G(n_195), .Q(n_25));
   DLH_X1 \Index_reg[6]  (.D(Index[6]), .G(n_195), .Q(n_26));
   DLH_X1 \Index_reg[5]  (.D(Index[5]), .G(n_195), .Q(n_27));
   DLH_X1 \Index_reg[4]  (.D(Index[4]), .G(n_195), .Q(n_28));
   DLH_X1 \Index_reg[3]  (.D(Index[3]), .G(n_195), .Q(n_29));
   DLH_X1 \Index_reg[2]  (.D(Index[2]), .G(n_195), .Q(n_30));
   DLH_X1 \Index_reg[1]  (.D(Index[1]), .G(n_195), .Q(n_31));
   DLH_X1 \Index_reg[0]  (.D(Index[0]), .G(n_195), .Q(n_32));
   datapath__0_59 i_29 (.Index({n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, 
      n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, 
      n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32}), 
      .p_0({n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, 
      n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, 
      n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33}));
   DLH_X1 \QuotientVar_reg[15]  (.D(QuotientVar[15]), .G(n_173), .Q(n_65));
   DLH_X1 \QuotientVar_reg[14]  (.D(QuotientVar[14]), .G(n_172), .Q(n_66));
   DLH_X1 \QuotientVar_reg[13]  (.D(QuotientVar[13]), .G(n_171), .Q(n_67));
   DLH_X1 \QuotientVar_reg[12]  (.D(QuotientVar[12]), .G(n_170), .Q(n_68));
   DLH_X1 \QuotientVar_reg[11]  (.D(QuotientVar[11]), .G(n_169), .Q(n_69));
   DLH_X1 \QuotientVar_reg[10]  (.D(QuotientVar[10]), .G(n_168), .Q(n_70));
   DLH_X1 \QuotientVar_reg[9]  (.D(QuotientVar[9]), .G(n_167), .Q(n_71));
   DLH_X1 \QuotientVar_reg[8]  (.D(QuotientVar[8]), .G(n_166), .Q(n_72));
   DLH_X1 \QuotientVar_reg[7]  (.D(QuotientVar[7]), .G(n_165), .Q(n_73));
   DLH_X1 \QuotientVar_reg[6]  (.D(QuotientVar[6]), .G(n_164), .Q(n_74));
   DLH_X1 \QuotientVar_reg[5]  (.D(QuotientVar[5]), .G(n_163), .Q(n_75));
   DLH_X1 \QuotientVar_reg[4]  (.D(QuotientVar[4]), .G(n_162), .Q(n_76));
   DLH_X1 \QuotientVar_reg[3]  (.D(QuotientVar[3]), .G(n_161), .Q(n_77));
   DLH_X1 \QuotientVar_reg[2]  (.D(QuotientVar[2]), .G(n_160), .Q(n_78));
   DLH_X1 \QuotientVar_reg[1]  (.D(QuotientVar[1]), .G(n_159), .Q(n_79));
   DLH_X1 \QuotientVar_reg[0]  (.D(QuotientVar[0]), .G(n_158), .Q(n_80));
   DLH_X1 \Divisor2_reg[28]  (.D(n_157), .G(n_195), .Q(n_81));
   DLH_X1 \Divisor2_reg[27]  (.D(n_156), .G(n_195), .Q(n_82));
   DLH_X1 \Divisor2_reg[26]  (.D(n_155), .G(n_195), .Q(n_83));
   DLH_X1 \Divisor2_reg[25]  (.D(n_154), .G(n_195), .Q(n_84));
   DLH_X1 \Divisor2_reg[24]  (.D(n_153), .G(n_195), .Q(n_85));
   DLH_X1 \Divisor2_reg[23]  (.D(n_152), .G(n_195), .Q(n_86));
   DLH_X1 \Divisor2_reg[22]  (.D(n_151), .G(n_195), .Q(n_87));
   DLH_X1 \Divisor2_reg[21]  (.D(n_150), .G(n_195), .Q(n_88));
   DLH_X1 \Divisor2_reg[20]  (.D(n_149), .G(n_195), .Q(n_89));
   DLH_X1 \Divisor2_reg[19]  (.D(n_148), .G(n_195), .Q(n_90));
   DLH_X1 \Divisor2_reg[18]  (.D(n_147), .G(n_195), .Q(n_91));
   DLH_X1 \Divisor2_reg[17]  (.D(n_146), .G(n_195), .Q(n_92));
   DLH_X1 \Divisor2_reg[16]  (.D(n_145), .G(n_195), .Q(n_93));
   DLH_X1 \Divisor2_reg[15]  (.D(n_144), .G(n_195), .Q(n_94));
   DLH_X1 \Divisor2_reg[14]  (.D(n_143), .G(n_195), .Q(n_95));
   DLH_X1 \Divisor2_reg[13]  (.D(n_142), .G(n_195), .Q(n_96));
   DLH_X1 \Divisor2_reg[12]  (.D(n_141), .G(n_195), .Q(n_97));
   DLH_X1 \Divisor2_reg[11]  (.D(n_140), .G(n_195), .Q(n_98));
   DLH_X1 \Divisor2_reg[10]  (.D(n_139), .G(n_195), .Q(n_99));
   DLH_X1 \Divisor2_reg[9]  (.D(n_138), .G(n_195), .Q(n_100));
   DLH_X1 \Divisor2_reg[8]  (.D(n_137), .G(n_195), .Q(n_101));
   DLH_X1 \Divisor2_reg[7]  (.D(n_136), .G(n_195), .Q(n_102));
   DLH_X1 \Divisor2_reg[6]  (.D(n_135), .G(n_195), .Q(n_103));
   DLH_X1 \Divisor2_reg[5]  (.D(n_134), .G(n_195), .Q(n_104));
   DLH_X1 \Divisor2_reg[4]  (.D(n_133), .G(n_195), .Q(n_105));
   DLH_X1 \Divisor2_reg[3]  (.D(n_132), .G(n_195), .Q(n_106));
   DLH_X1 \Divisor2_reg[2]  (.D(n_131), .G(n_195), .Q(n_107));
   DLH_X1 \Divisor2_reg[1]  (.D(n_130), .G(n_195), .Q(n_108));
   DLH_X1 \Divisor2_reg[0]  (.D(n_129), .G(n_195), .Q(n_109));
   DLH_X1 \Dividend2_reg[15]  (.D(Dividend2[15]), .G(n_128), .Q(n_110));
   DLH_X1 \Dividend2_reg[14]  (.D(Dividend2[14]), .G(n_128), .Q(n_111));
   DLH_X1 \Dividend2_reg[13]  (.D(Dividend2[13]), .G(n_128), .Q(n_112));
   DLH_X1 \Dividend2_reg[12]  (.D(Dividend2[12]), .G(n_128), .Q(n_113));
   DLH_X1 \Dividend2_reg[11]  (.D(Dividend2[11]), .G(n_128), .Q(n_114));
   DLH_X1 \Dividend2_reg[10]  (.D(Dividend2[10]), .G(n_128), .Q(n_115));
   DLH_X1 \Dividend2_reg[9]  (.D(Dividend2[9]), .G(n_128), .Q(n_116));
   DLH_X1 \Dividend2_reg[8]  (.D(Dividend2[8]), .G(n_128), .Q(n_117));
   DLH_X1 \Dividend2_reg[7]  (.D(Dividend2[7]), .G(n_128), .Q(n_118));
   DLH_X1 \Dividend2_reg[6]  (.D(Dividend2[6]), .G(n_128), .Q(n_119));
   DLH_X1 \Dividend2_reg[5]  (.D(Dividend2[5]), .G(n_128), .Q(n_120));
   DLH_X1 \Dividend2_reg[4]  (.D(Dividend2[4]), .G(n_128), .Q(n_121));
   DLH_X1 \Dividend2_reg[3]  (.D(Dividend2[3]), .G(n_128), .Q(n_122));
   DLH_X1 \Dividend2_reg[2]  (.D(Dividend2[2]), .G(n_128), .Q(n_123));
   DLH_X1 \Dividend2_reg[1]  (.D(Dividend2[1]), .G(n_128), .Q(n_124));
   DLH_X1 \Dividend2_reg[0]  (.D(Dividend2[0]), .G(n_128), .Q(n_125));
   DLH_X1 FIRST_ONE_reg (.D(FIRST_ONE), .G(n_127), .Q(n_126));
   HA_X1 i_0_0 (.A(n_0_13), .B(n_0_14__0), .CO(n_0_19__0), .S());
   FA_X1 i_0_1 (.A(n_0_15), .B(n_0_16), .CI(n_0_19__0), .CO(n_0_20), .S());
   HA_X1 i_0_2 (.A(n_0_26), .B(n_0_10), .CO(n_0_0), .S());
   HA_X1 i_0_3 (.A(n_0_7), .B(n_0_0), .CO(n_0_1), .S());
   NAND2_X1 i_0_4 (.A1(n_0_2), .A2(n_0_245), .ZN(n_0_16));
   XNOR2_X1 i_0_5 (.A(n_0_253), .B(n_0_110), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(n_0_15), .A2(n_0_3), .ZN(n_0_14__0));
   NAND2_X1 i_0_7 (.A1(n_0_5), .A2(n_0_4__0), .ZN(n_0_3));
   OR2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_4__0), .ZN(n_0_15));
   XNOR2_X1 i_0_9 (.A(n_0_253), .B(n_0_245), .ZN(n_0_4__0));
   NAND4_X1 i_0_10 (.A1(n_0_25), .A2(n_0_9__0), .A3(n_0_6), .A4(n_0_5), .ZN(
      n_0_13));
   OR2_X1 i_0_11 (.A1(n_0_7), .A2(n_0_225), .ZN(n_0_5));
   NAND2_X1 i_0_12 (.A1(n_0_7), .A2(n_0_225), .ZN(n_0_6));
   OR3_X1 i_0_13 (.A1(Divisor[14]), .A2(n_0_8), .A3(n_0_246), .ZN(n_0_7));
   AOI21_X1 i_0_14 (.A(n_0_247), .B1(n_0_112), .B2(n_0_243), .ZN(n_0_8));
   OAI211_X1 i_0_15 (.A(n_0_232), .B(n_0_10), .C1(n_0_26), .C2(n_0_228), 
      .ZN(n_0_9__0));
   OAI21_X1 i_0_16 (.A(n_0_11), .B1(n_0_12), .B2(Divisor[14]), .ZN(n_0_10));
   OAI21_X1 i_0_17 (.A(n_0_245), .B1(n_0_21), .B2(Divisor[7]), .ZN(n_0_11));
   NOR2_X1 i_0_18 (.A1(Divisor[13]), .A2(n_0_17), .ZN(n_0_12));
   NOR2_X1 i_0_19 (.A1(Divisor[12]), .A2(n_0_18), .ZN(n_0_17));
   AOI21_X1 i_0_20 (.A(Divisor[11]), .B1(n_0_290), .B2(Divisor[9]), .ZN(n_0_18));
   NOR2_X1 i_0_21 (.A1(Divisor[6]), .A2(n_0_22), .ZN(n_0_21));
   NOR2_X1 i_0_22 (.A1(Divisor[5]), .A2(n_0_23), .ZN(n_0_22));
   NOR2_X1 i_0_23 (.A1(Divisor[4]), .A2(n_0_24__0), .ZN(n_0_23));
   AOI21_X1 i_0_24 (.A(Divisor[3]), .B1(n_0_289), .B2(Divisor[1]), .ZN(n_0_24__0));
   NAND2_X1 i_0_25 (.A1(n_0_26), .A2(n_0_228), .ZN(n_0_25));
   OAI21_X1 i_0_26 (.A(n_0_27), .B1(n_0_246), .B2(n_0_249), .ZN(n_0_26));
   AOI21_X1 i_0_27 (.A(Divisor[14]), .B1(n_0_28), .B2(n_0_245), .ZN(n_0_27));
   OR3_X1 i_0_28 (.A1(Divisor[7]), .A2(Divisor[6]), .A3(n_0_29__0), .ZN(n_0_28));
   NOR3_X1 i_0_29 (.A1(Divisor[5]), .A2(Divisor[4]), .A3(n_0_244), .ZN(n_0_29__0));
   NOR3_X1 i_0_30 (.A1(Reset), .A2(n_0_203), .A3(n_0_30), .ZN(n_127));
   NOR3_X1 i_0_31 (.A1(n_0), .A2(n_126), .A3(n_0_161), .ZN(n_0_30));
   AOI21_X1 i_0_32 (.A(Reset), .B1(n_0_105), .B2(n_0_31), .ZN(n_128));
   NAND2_X1 i_0_33 (.A1(n_0_286), .A2(n_126), .ZN(n_0_31));
   OAI21_X1 i_0_34 (.A(n_0_128), .B1(n_0_278), .B2(n_0), .ZN(Dividend2[0]));
   OAI21_X1 i_0_35 (.A(n_0_34__0), .B1(n_0_32), .B2(n_0_313), .ZN(Dividend2[1]));
   XNOR2_X1 i_0_36 (.A(n_0_293), .B(n_0_33), .ZN(n_0_32));
   NAND2_X1 i_0_37 (.A1(Dividend[15]), .A2(Dividend[0]), .ZN(n_0_33));
   NAND2_X1 i_0_38 (.A1(n_0_286), .A2(addOut[1]), .ZN(n_0_34__0));
   OAI21_X1 i_0_39 (.A(n_0_36), .B1(n_0_35), .B2(n_0_313), .ZN(Dividend2[2]));
   XNOR2_X1 i_0_40 (.A(n_0_294), .B(n_0_40), .ZN(n_0_35));
   NAND2_X1 i_0_41 (.A1(n_0_286), .A2(addOut[2]), .ZN(n_0_36));
   OAI21_X1 i_0_42 (.A(n_0_37), .B1(n_0_38), .B2(n_0_313), .ZN(Dividend2[3]));
   NAND2_X1 i_0_43 (.A1(n_0_286), .A2(addOut[3]), .ZN(n_0_37));
   XNOR2_X1 i_0_44 (.A(Dividend[3]), .B(n_0_39__0), .ZN(n_0_38));
   OAI21_X1 i_0_45 (.A(n_0_40), .B1(n_0_294), .B2(n_0_307), .ZN(n_0_39__0));
   OAI21_X1 i_0_46 (.A(Dividend[15]), .B1(Dividend[1]), .B2(Dividend[0]), 
      .ZN(n_0_40));
   OAI22_X1 i_0_47 (.A1(n_0_313), .A2(n_0_41), .B1(n_0), .B2(n_0_279), .ZN(
      Dividend2[4]));
   XNOR2_X1 i_0_48 (.A(n_0_296), .B(n_0_44__0), .ZN(n_0_41));
   OAI22_X1 i_0_49 (.A1(n_0_313), .A2(n_0_42), .B1(n_0), .B2(n_0_280), .ZN(
      Dividend2[5]));
   XNOR2_X1 i_0_50 (.A(n_0_297), .B(n_0_43), .ZN(n_0_42));
   OAI21_X1 i_0_51 (.A(Dividend[15]), .B1(n_0_261), .B2(Dividend[4]), .ZN(n_0_43));
   NAND2_X1 i_0_52 (.A1(n_0_261), .A2(Dividend[15]), .ZN(n_0_44__0));
   OAI21_X1 i_0_53 (.A(n_0_46), .B1(n_0_45), .B2(n_0_313), .ZN(Dividend2[6]));
   XNOR2_X1 i_0_54 (.A(n_0_298), .B(n_0_50), .ZN(n_0_45));
   NAND2_X1 i_0_55 (.A1(n_0_286), .A2(addOut[6]), .ZN(n_0_46));
   OAI21_X1 i_0_56 (.A(n_0_48), .B1(n_0_47), .B2(n_0_313), .ZN(Dividend2[7]));
   XNOR2_X1 i_0_57 (.A(n_0_299), .B(n_0_49__0), .ZN(n_0_47));
   NAND2_X1 i_0_58 (.A1(n_0_286), .A2(addOut[7]), .ZN(n_0_48));
   OAI21_X1 i_0_59 (.A(Dividend[15]), .B1(n_0_259), .B2(Dividend[6]), .ZN(
      n_0_49__0));
   NAND2_X1 i_0_60 (.A1(n_0_259), .A2(Dividend[15]), .ZN(n_0_50));
   OAI22_X1 i_0_61 (.A1(n_0_313), .A2(n_0_51), .B1(n_0), .B2(n_0_281), .ZN(
      Dividend2[8]));
   XNOR2_X1 i_0_62 (.A(n_0_300), .B(n_0_68), .ZN(n_0_51));
   OAI22_X1 i_0_63 (.A1(n_0_313), .A2(n_0_52), .B1(n_0), .B2(n_0_282), .ZN(
      Dividend2[9]));
   XNOR2_X1 i_0_64 (.A(n_0_301), .B(n_0_53), .ZN(n_0_52));
   OAI21_X1 i_0_65 (.A(Dividend[15]), .B1(n_0_257), .B2(Dividend[8]), .ZN(n_0_53));
   OAI21_X1 i_0_66 (.A(n_0_55), .B1(n_0_54__0), .B2(n_0_313), .ZN(Dividend2[10]));
   XNOR2_X1 i_0_67 (.A(n_0_302), .B(n_0_59__0), .ZN(n_0_54__0));
   NAND2_X1 i_0_68 (.A1(n_0_286), .A2(addOut[10]), .ZN(n_0_55));
   OAI21_X1 i_0_69 (.A(n_0_57), .B1(n_0_56), .B2(n_0_313), .ZN(Dividend2[11]));
   XNOR2_X1 i_0_70 (.A(n_0_303), .B(n_0_58), .ZN(n_0_56));
   NAND2_X1 i_0_71 (.A1(n_0_286), .A2(addOut[11]), .ZN(n_0_57));
   OAI21_X1 i_0_72 (.A(Dividend[15]), .B1(n_0_252), .B2(Dividend[10]), .ZN(
      n_0_58));
   NAND2_X1 i_0_73 (.A1(n_0_252), .A2(Dividend[15]), .ZN(n_0_59__0));
   OAI22_X1 i_0_74 (.A1(n_0_313), .A2(n_0_60), .B1(n_0), .B2(n_0_283), .ZN(
      Dividend2[12]));
   XNOR2_X1 i_0_75 (.A(n_0_304), .B(n_0_67), .ZN(n_0_60));
   OAI21_X1 i_0_76 (.A(n_0_62), .B1(n_0_61), .B2(n_0_313), .ZN(Dividend2[13]));
   XNOR2_X1 i_0_77 (.A(n_0_305), .B(n_0_63), .ZN(n_0_61));
   NAND2_X1 i_0_78 (.A1(n_0_286), .A2(addOut[13]), .ZN(n_0_62));
   OAI21_X1 i_0_79 (.A(Dividend[15]), .B1(n_0_251), .B2(Dividend[12]), .ZN(
      n_0_63));
   OAI21_X1 i_0_80 (.A(n_0_65), .B1(n_0_64__0), .B2(n_0_313), .ZN(Dividend2[14]));
   XNOR2_X1 i_0_81 (.A(Dividend[14]), .B(n_0_66), .ZN(n_0_64__0));
   NAND2_X1 i_0_82 (.A1(n_0_286), .A2(addOut[14]), .ZN(n_0_65));
   OAI21_X1 i_0_83 (.A(n_0_67), .B1(n_0_256), .B2(n_0_307), .ZN(n_0_66));
   NAND2_X1 i_0_84 (.A1(n_0_251), .A2(Dividend[15]), .ZN(n_0_67));
   NAND2_X1 i_0_85 (.A1(n_0_257), .A2(Dividend[15]), .ZN(n_0_68));
   OAI21_X1 i_0_86 (.A(n_0_69__0), .B1(n_0_284), .B2(n_0), .ZN(Dividend2[15]));
   NAND3_X1 i_0_87 (.A1(Dividend[15]), .A2(n_0_262), .A3(n_0_250), .ZN(n_0_69__0));
   NOR2_X1 i_0_88 (.A1(n_0_4__1), .A2(n_0), .ZN(n_129));
   NOR2_X1 i_0_89 (.A1(n_0_9__1), .A2(n_0), .ZN(n_130));
   NOR2_X1 i_0_90 (.A1(n_0_14__1), .A2(n_0), .ZN(n_131));
   NOR2_X1 i_0_91 (.A1(n_0_19__1), .A2(n_0), .ZN(n_132));
   NOR2_X1 i_0_92 (.A1(n_0_24__1), .A2(n_0), .ZN(n_133));
   NOR2_X1 i_0_93 (.A1(n_0_29__1), .A2(n_0), .ZN(n_134));
   NOR2_X1 i_0_94 (.A1(n_0_34__1), .A2(n_0), .ZN(n_135));
   NOR2_X1 i_0_95 (.A1(n_0_39__1), .A2(n_0), .ZN(n_136));
   NOR2_X1 i_0_96 (.A1(n_0_44__1), .A2(n_0), .ZN(n_137));
   NOR2_X1 i_0_97 (.A1(n_0_49__1), .A2(n_0), .ZN(n_138));
   NOR2_X1 i_0_98 (.A1(n_0_54__1), .A2(n_0), .ZN(n_139));
   NOR2_X1 i_0_99 (.A1(n_0_59__1), .A2(n_0), .ZN(n_140));
   NOR2_X1 i_0_100 (.A1(n_0_64__1), .A2(n_0), .ZN(n_141));
   NOR2_X1 i_0_101 (.A1(n_0_69__1), .A2(n_0), .ZN(n_142));
   OAI22_X1 i_0_102 (.A1(n_0_287), .A2(n_0_105), .B1(n_0), .B2(n_0_74__1), 
      .ZN(n_143));
   OAI21_X1 i_0_103 (.A(n_0_72), .B1(n_0_105), .B2(n_0_70), .ZN(n_144));
   XNOR2_X1 i_0_104 (.A(n_0_288), .B(n_0_71), .ZN(n_0_70));
   NAND2_X1 i_0_105 (.A1(Divisor[15]), .A2(Divisor[0]), .ZN(n_0_71));
   NAND2_X1 i_0_106 (.A1(n_0_286), .A2(n_93), .ZN(n_0_72));
   OAI22_X1 i_0_107 (.A1(n_0_105), .A2(n_0_73), .B1(n_0_309), .B2(n_0), .ZN(
      n_145));
   XNOR2_X1 i_0_108 (.A(n_0_289), .B(n_0_76), .ZN(n_0_73));
   OAI22_X1 i_0_109 (.A1(n_0_105), .A2(n_0_74__0), .B1(n_0_310), .B2(n_0), 
      .ZN(n_146));
   XNOR2_X1 i_0_110 (.A(Divisor[3]), .B(n_0_75), .ZN(n_0_74__0));
   OAI21_X1 i_0_111 (.A(n_0_76), .B1(n_0_289), .B2(n_0_291), .ZN(n_0_75));
   OAI21_X1 i_0_112 (.A(Divisor[15]), .B1(Divisor[1]), .B2(Divisor[0]), .ZN(
      n_0_76));
   OAI21_X1 i_0_113 (.A(n_0_78), .B1(n_0_105), .B2(n_0_77), .ZN(n_147));
   XOR2_X1 i_0_114 (.A(Divisor[4]), .B(n_0_81), .Z(n_0_77));
   NAND2_X1 i_0_115 (.A1(n_0_286), .A2(n_90), .ZN(n_0_78));
   OAI22_X1 i_0_116 (.A1(n_0_105), .A2(n_0_79), .B1(n_0_311), .B2(n_0), .ZN(
      n_148));
   XOR2_X1 i_0_117 (.A(Divisor[5]), .B(n_0_80), .Z(n_0_79));
   OAI21_X1 i_0_118 (.A(Divisor[15]), .B1(n_0_243), .B2(Divisor[4]), .ZN(n_0_80));
   NAND2_X1 i_0_119 (.A1(n_0_243), .A2(Divisor[15]), .ZN(n_0_81));
   OAI22_X1 i_0_120 (.A1(n_0_105), .A2(n_0_82), .B1(n_0_312), .B2(n_0), .ZN(
      n_149));
   XOR2_X1 i_0_121 (.A(Divisor[6]), .B(n_0_83), .Z(n_0_82));
   NAND2_X1 i_0_122 (.A1(n_0_242), .A2(Divisor[15]), .ZN(n_0_83));
   OAI21_X1 i_0_123 (.A(n_0_86), .B1(n_0_84), .B2(n_0_105), .ZN(n_150));
   XOR2_X1 i_0_124 (.A(Divisor[7]), .B(n_0_85), .Z(n_0_84));
   NAND2_X1 i_0_125 (.A1(n_0_241), .A2(Divisor[15]), .ZN(n_0_85));
   NAND2_X1 i_0_126 (.A1(n_0_286), .A2(n_87), .ZN(n_0_86));
   OAI21_X1 i_0_127 (.A(n_0_88), .B1(n_0_87), .B2(n_0_105), .ZN(n_151));
   XNOR2_X1 i_0_128 (.A(Divisor[8]), .B(n_0_97), .ZN(n_0_87));
   NAND2_X1 i_0_129 (.A1(n_0_286), .A2(n_86), .ZN(n_0_88));
   OAI21_X1 i_0_130 (.A(n_0_90), .B1(n_0_89), .B2(n_0_105), .ZN(n_152));
   XOR2_X1 i_0_131 (.A(Divisor[9]), .B(n_0_96), .Z(n_0_89));
   NAND2_X1 i_0_132 (.A1(n_0_286), .A2(n_85), .ZN(n_0_90));
   OAI21_X1 i_0_133 (.A(n_0_92), .B1(n_0_91), .B2(n_0_105), .ZN(n_153));
   XNOR2_X1 i_0_134 (.A(n_0_290), .B(n_0_95), .ZN(n_0_91));
   NAND2_X1 i_0_135 (.A1(n_0_286), .A2(n_84), .ZN(n_0_92));
   OAI21_X1 i_0_136 (.A(n_0_98), .B1(n_0_93), .B2(n_0_105), .ZN(n_154));
   XOR2_X1 i_0_137 (.A(Divisor[11]), .B(n_0_94), .Z(n_0_93));
   OAI21_X1 i_0_138 (.A(Divisor[15]), .B1(n_0_109), .B2(Divisor[10]), .ZN(n_0_94));
   NAND2_X1 i_0_139 (.A1(n_0_109), .A2(Divisor[15]), .ZN(n_0_95));
   OAI21_X1 i_0_140 (.A(Divisor[15]), .B1(n_0_110), .B2(Divisor[8]), .ZN(n_0_96));
   NOR2_X1 i_0_141 (.A1(n_0_111), .A2(n_0_291), .ZN(n_0_97));
   NAND2_X1 i_0_142 (.A1(n_0_286), .A2(n_83), .ZN(n_0_98));
   OAI21_X1 i_0_143 (.A(n_0_100), .B1(n_0_99), .B2(n_0_105), .ZN(n_155));
   XOR2_X1 i_0_144 (.A(Divisor[12]), .B(n_0_107), .Z(n_0_99));
   NAND2_X1 i_0_145 (.A1(n_0_286), .A2(n_82), .ZN(n_0_100));
   OAI21_X1 i_0_146 (.A(n_0_103), .B1(n_0_101), .B2(n_0_105), .ZN(n_156));
   XOR2_X1 i_0_147 (.A(Divisor[13]), .B(n_0_102), .Z(n_0_101));
   OAI21_X1 i_0_148 (.A(Divisor[15]), .B1(n_0_108), .B2(Divisor[12]), .ZN(
      n_0_102));
   NAND2_X1 i_0_149 (.A1(n_0_286), .A2(n_81), .ZN(n_0_103));
   NOR2_X1 i_0_150 (.A1(n_0_105), .A2(n_0_104), .ZN(n_157));
   XOR2_X1 i_0_151 (.A(Divisor[14]), .B(n_0_106), .Z(n_0_104));
   NAND2_X1 i_0_152 (.A1(n_0_262), .A2(n_0_239), .ZN(n_0_105));
   OAI21_X1 i_0_153 (.A(Divisor[15]), .B1(n_0_246), .B2(n_0_108), .ZN(n_0_106));
   NAND2_X1 i_0_154 (.A1(n_0_108), .A2(Divisor[15]), .ZN(n_0_107));
   NAND3_X1 i_0_155 (.A1(n_0_249), .A2(n_0_248), .A3(n_0_111), .ZN(n_0_108));
   NAND2_X1 i_0_156 (.A1(n_0_248), .A2(n_0_111), .ZN(n_0_109));
   INV_X1 i_0_157 (.A(n_0_111), .ZN(n_0_110));
   NOR2_X1 i_0_158 (.A1(n_0_241), .A2(Divisor[7]), .ZN(n_0_111));
   NOR4_X1 i_0_159 (.A1(Divisor[7]), .A2(Divisor[6]), .A3(Divisor[5]), .A4(
      Divisor[4]), .ZN(n_0_112));
   OAI21_X1 i_0_160 (.A(n_0_122), .B1(n_0_115), .B2(n_0_206), .ZN(n_158));
   OAI21_X1 i_0_161 (.A(n_0_122), .B1(n_0_116), .B2(n_0_206), .ZN(n_159));
   OAI21_X1 i_0_162 (.A(n_0_122), .B1(n_0_118), .B2(n_0_206), .ZN(n_160));
   OAI21_X1 i_0_163 (.A(n_0_122), .B1(n_0_119), .B2(n_0_206), .ZN(n_161));
   OAI21_X1 i_0_164 (.A(n_0_122), .B1(n_0_115), .B2(n_0_113), .ZN(n_162));
   OAI21_X1 i_0_165 (.A(n_0_122), .B1(n_0_116), .B2(n_0_113), .ZN(n_163));
   OAI21_X1 i_0_166 (.A(n_0_122), .B1(n_0_118), .B2(n_0_113), .ZN(n_164));
   OAI21_X1 i_0_167 (.A(n_0_122), .B1(n_0_119), .B2(n_0_113), .ZN(n_165));
   OR3_X1 i_0_168 (.A1(n_0_207), .A2(n_29), .A3(n_0_308), .ZN(n_0_113));
   OAI21_X1 i_0_169 (.A(n_0_122), .B1(n_0_115), .B2(n_0_114), .ZN(n_166));
   OAI21_X1 i_0_170 (.A(n_0_122), .B1(n_0_116), .B2(n_0_114), .ZN(n_167));
   OAI21_X1 i_0_171 (.A(n_0_122), .B1(n_0_118), .B2(n_0_114), .ZN(n_168));
   OAI21_X1 i_0_172 (.A(n_0_122), .B1(n_0_119), .B2(n_0_114), .ZN(n_169));
   NAND3_X1 i_0_173 (.A1(n_29), .A2(n_0_208), .A3(n_0_308), .ZN(n_0_114));
   OAI21_X1 i_0_174 (.A(n_0_122), .B1(n_0_121), .B2(n_0_115), .ZN(n_170));
   NAND2_X1 i_0_175 (.A1(n_33), .A2(n_0_117), .ZN(n_0_115));
   OAI21_X1 i_0_176 (.A(n_0_122), .B1(n_0_121), .B2(n_0_116), .ZN(n_171));
   NAND2_X1 i_0_177 (.A1(n_32), .A2(n_0_117), .ZN(n_0_116));
   NOR2_X1 i_0_178 (.A1(n_0_123), .A2(n_31), .ZN(n_0_117));
   OAI21_X1 i_0_179 (.A(n_0_122), .B1(n_0_121), .B2(n_0_118), .ZN(n_172));
   NAND2_X1 i_0_180 (.A1(n_33), .A2(n_0_120), .ZN(n_0_118));
   OAI21_X1 i_0_181 (.A(n_0_122), .B1(n_0_121), .B2(n_0_119), .ZN(n_173));
   NAND2_X1 i_0_182 (.A1(n_32), .A2(n_0_120), .ZN(n_0_119));
   AND2_X1 i_0_183 (.A1(n_31), .A2(n_176), .ZN(n_0_120));
   NAND3_X1 i_0_184 (.A1(n_29), .A2(n_30), .A3(n_0_208), .ZN(n_0_121));
   NAND2_X1 i_0_185 (.A1(n_0_262), .A2(n_0_285), .ZN(n_0_122));
   OAI21_X1 i_0_186 (.A(n_0), .B1(n_0_125), .B2(n_0_292), .ZN(QuotientVar[0]));
   OAI21_X1 i_0_187 (.A(n_0), .B1(n_0_125), .B2(n_0_293), .ZN(QuotientVar[1]));
   OAI21_X1 i_0_188 (.A(n_0), .B1(n_0_125), .B2(n_0_294), .ZN(QuotientVar[2]));
   OAI21_X1 i_0_189 (.A(n_0), .B1(n_0_125), .B2(n_0_295), .ZN(QuotientVar[3]));
   OAI21_X1 i_0_190 (.A(n_0), .B1(n_0_125), .B2(n_0_296), .ZN(QuotientVar[4]));
   OAI21_X1 i_0_191 (.A(n_0), .B1(n_0_125), .B2(n_0_297), .ZN(QuotientVar[5]));
   OAI21_X1 i_0_192 (.A(n_0), .B1(n_0_125), .B2(n_0_298), .ZN(QuotientVar[6]));
   OAI21_X1 i_0_193 (.A(n_0), .B1(n_0_125), .B2(n_0_299), .ZN(QuotientVar[7]));
   OAI21_X1 i_0_194 (.A(n_0), .B1(n_0_125), .B2(n_0_300), .ZN(QuotientVar[8]));
   OAI21_X1 i_0_195 (.A(n_0), .B1(n_0_125), .B2(n_0_301), .ZN(QuotientVar[9]));
   OAI21_X1 i_0_196 (.A(n_0), .B1(n_0_125), .B2(n_0_302), .ZN(QuotientVar[10]));
   OAI21_X1 i_0_197 (.A(n_0), .B1(n_0_125), .B2(n_0_303), .ZN(QuotientVar[11]));
   OAI21_X1 i_0_198 (.A(n_0), .B1(n_0_125), .B2(n_0_304), .ZN(QuotientVar[12]));
   OAI21_X1 i_0_199 (.A(n_0), .B1(n_0_125), .B2(n_0_305), .ZN(QuotientVar[13]));
   OAI21_X1 i_0_200 (.A(n_0), .B1(n_0_125), .B2(n_0_306), .ZN(QuotientVar[14]));
   OAI21_X1 i_0_201 (.A(n_0_313), .B1(n_0), .B2(n_32), .ZN(Index[0]));
   AND2_X1 i_0_202 (.A1(n_0_286), .A2(n_34), .ZN(Index[1]));
   OAI21_X1 i_0_203 (.A(n_0_313), .B1(n_0_271), .B2(n_0), .ZN(Index[2]));
   AND2_X1 i_0_204 (.A1(n_0_286), .A2(n_36), .ZN(Index[3]));
   OAI21_X1 i_0_205 (.A(n_0_313), .B1(n_0_272), .B2(n_0), .ZN(Index[4]));
   AND2_X1 i_0_206 (.A1(n_0_286), .A2(n_38), .ZN(Index[5]));
   AND2_X1 i_0_207 (.A1(n_0_286), .A2(n_39), .ZN(Index[6]));
   AND2_X1 i_0_208 (.A1(n_0_286), .A2(n_40), .ZN(Index[7]));
   AND2_X1 i_0_209 (.A1(n_0_286), .A2(n_41), .ZN(Index[8]));
   AND2_X1 i_0_210 (.A1(n_0_286), .A2(n_42), .ZN(Index[9]));
   AND2_X1 i_0_211 (.A1(n_0_286), .A2(n_43), .ZN(Index[10]));
   AND2_X1 i_0_212 (.A1(n_0_286), .A2(n_44), .ZN(Index[11]));
   AND2_X1 i_0_213 (.A1(n_0_286), .A2(n_45), .ZN(Index[12]));
   AND2_X1 i_0_214 (.A1(n_0_286), .A2(n_46), .ZN(Index[13]));
   AND2_X1 i_0_215 (.A1(n_0_286), .A2(n_47), .ZN(Index[14]));
   AND2_X1 i_0_216 (.A1(n_0_286), .A2(n_48), .ZN(Index[15]));
   AND2_X1 i_0_217 (.A1(n_0_286), .A2(n_49), .ZN(Index[16]));
   AND2_X1 i_0_218 (.A1(n_0_286), .A2(n_50), .ZN(Index[17]));
   AND2_X1 i_0_219 (.A1(n_0_286), .A2(n_51), .ZN(Index[18]));
   AND2_X1 i_0_220 (.A1(n_0_286), .A2(n_52), .ZN(Index[19]));
   AND2_X1 i_0_221 (.A1(n_0_286), .A2(n_53), .ZN(Index[20]));
   AND2_X1 i_0_222 (.A1(n_0_286), .A2(n_54), .ZN(Index[21]));
   AND2_X1 i_0_223 (.A1(n_0_286), .A2(n_55), .ZN(Index[22]));
   AND2_X1 i_0_224 (.A1(n_0_286), .A2(n_56), .ZN(Index[23]));
   AND2_X1 i_0_225 (.A1(n_0_286), .A2(n_57), .ZN(Index[24]));
   AND2_X1 i_0_226 (.A1(n_0_286), .A2(n_58), .ZN(Index[25]));
   AND2_X1 i_0_227 (.A1(n_0_286), .A2(n_59), .ZN(Index[26]));
   AND2_X1 i_0_228 (.A1(n_0_286), .A2(n_60), .ZN(Index[27]));
   AND2_X1 i_0_229 (.A1(n_0_286), .A2(n_61), .ZN(Index[28]));
   AND2_X1 i_0_230 (.A1(n_0_286), .A2(n_62), .ZN(Index[29]));
   AND2_X1 i_0_231 (.A1(n_0_286), .A2(n_63), .ZN(Index[30]));
   AND2_X1 i_0_232 (.A1(n_0_286), .A2(n_64), .ZN(Index[31]));
   NAND2_X1 i_0_233 (.A1(n_0_203), .A2(n_0_285), .ZN(n_174));
   OAI211_X1 i_0_234 (.A(n_0_285), .B(n_0_204), .C1(n_0_222), .C2(n_0_313), 
      .ZN(n_175));
   INV_X1 i_0_235 (.A(n_0_123), .ZN(n_176));
   NAND2_X1 i_0_236 (.A1(FIRST_ONE), .A2(n_0_285), .ZN(n_0_123));
   INV_X1 i_0_237 (.A(n_0_124), .ZN(FIRST_ONE));
   NAND2_X1 i_0_238 (.A1(n_0_161), .A2(n_0_286), .ZN(n_0_124));
   AOI21_X1 i_0_239 (.A(Reset), .B1(n_0_204), .B2(n_0_125), .ZN(n_177));
   OAI21_X1 i_0_240 (.A(n_0_262), .B1(n_0_250), .B2(n_0_126), .ZN(n_0_125));
   NOR3_X1 i_0_241 (.A1(n_0_241), .A2(n_0_127), .A3(Divisor[15]), .ZN(n_0_126));
   NAND2_X1 i_0_242 (.A1(Divisor[7]), .A2(n_0_245), .ZN(n_0_127));
   OAI21_X1 i_0_243 (.A(n_0_128), .B1(n_0_160), .B2(n_0), .ZN(n_178));
   NAND2_X1 i_0_244 (.A1(Dividend[0]), .A2(n_0_262), .ZN(n_0_128));
   OAI22_X1 i_0_245 (.A1(n_0_129), .A2(n_0), .B1(n_0_293), .B2(n_0_313), 
      .ZN(n_179));
   XNOR2_X1 i_0_246 (.A(n_79), .B(n_0_159), .ZN(n_0_129));
   OAI22_X1 i_0_247 (.A1(n_0_130), .A2(n_0), .B1(n_0_294), .B2(n_0_313), 
      .ZN(n_180));
   XOR2_X1 i_0_248 (.A(n_78), .B(n_0_158), .Z(n_0_130));
   OAI22_X1 i_0_249 (.A1(n_0_131), .A2(n_0), .B1(n_0_295), .B2(n_0_313), 
      .ZN(n_181));
   XOR2_X1 i_0_250 (.A(n_77), .B(n_0_156), .Z(n_0_131));
   OAI22_X1 i_0_251 (.A1(n_0_132), .A2(n_0), .B1(n_0_296), .B2(n_0_313), 
      .ZN(n_182));
   XNOR2_X1 i_0_252 (.A(n_76), .B(n_0_155), .ZN(n_0_132));
   OAI22_X1 i_0_253 (.A1(n_0_133), .A2(n_0), .B1(n_0_297), .B2(n_0_313), 
      .ZN(n_183));
   XNOR2_X1 i_0_254 (.A(n_75), .B(n_0_154), .ZN(n_0_133));
   OAI22_X1 i_0_255 (.A1(n_0_134), .A2(n_0), .B1(n_0_298), .B2(n_0_313), 
      .ZN(n_184));
   XNOR2_X1 i_0_256 (.A(n_0_274), .B(n_0_153), .ZN(n_0_134));
   OAI22_X1 i_0_257 (.A1(n_0_135), .A2(n_0), .B1(n_0_299), .B2(n_0_313), 
      .ZN(n_185));
   XNOR2_X1 i_0_258 (.A(n_73), .B(n_0_152), .ZN(n_0_135));
   OAI22_X1 i_0_259 (.A1(n_0_136), .A2(n_0), .B1(n_0_300), .B2(n_0_313), 
      .ZN(n_186));
   XNOR2_X1 i_0_260 (.A(n_72), .B(n_0_150), .ZN(n_0_136));
   OAI22_X1 i_0_261 (.A1(n_0_137), .A2(n_0), .B1(n_0_301), .B2(n_0_313), 
      .ZN(n_187));
   XNOR2_X1 i_0_262 (.A(n_0_275), .B(n_0_149), .ZN(n_0_137));
   OAI22_X1 i_0_263 (.A1(n_0_138), .A2(n_0), .B1(n_0_302), .B2(n_0_313), 
      .ZN(n_188));
   XNOR2_X1 i_0_264 (.A(n_70), .B(n_0_148), .ZN(n_0_138));
   OAI22_X1 i_0_265 (.A1(n_0_139), .A2(n_0), .B1(n_0_303), .B2(n_0_313), 
      .ZN(n_189));
   XNOR2_X1 i_0_266 (.A(n_69), .B(n_0_146), .ZN(n_0_139));
   OAI22_X1 i_0_267 (.A1(n_0_140), .A2(n_0), .B1(n_0_304), .B2(n_0_313), 
      .ZN(n_190));
   XNOR2_X1 i_0_268 (.A(n_0_276), .B(n_0_145), .ZN(n_0_140));
   OAI22_X1 i_0_269 (.A1(n_0_141), .A2(n_0), .B1(n_0_305), .B2(n_0_313), 
      .ZN(n_191));
   XNOR2_X1 i_0_270 (.A(n_67), .B(n_0_144), .ZN(n_0_141));
   OAI22_X1 i_0_271 (.A1(n_0_142), .A2(n_0), .B1(n_0_306), .B2(n_0_313), 
      .ZN(n_192));
   XOR2_X1 i_0_272 (.A(n_66), .B(n_0_143), .Z(n_0_142));
   AOI21_X1 i_0_273 (.A(n_0_144), .B1(n_0_200), .B2(n_67), .ZN(n_0_143));
   OAI21_X1 i_0_274 (.A(n_0_145), .B1(n_0_199), .B2(n_0_276), .ZN(n_0_144));
   AOI21_X1 i_0_275 (.A(n_0_146), .B1(n_0_200), .B2(n_69), .ZN(n_0_145));
   INV_X1 i_0_276 (.A(n_0_147), .ZN(n_0_146));
   AOI21_X1 i_0_277 (.A(n_0_148), .B1(n_0_200), .B2(n_70), .ZN(n_0_147));
   OAI21_X1 i_0_278 (.A(n_0_149), .B1(n_0_199), .B2(n_0_275), .ZN(n_0_148));
   AOI21_X1 i_0_279 (.A(n_0_150), .B1(n_0_200), .B2(n_72), .ZN(n_0_149));
   INV_X1 i_0_280 (.A(n_0_151), .ZN(n_0_150));
   AOI21_X1 i_0_281 (.A(n_0_152), .B1(n_0_200), .B2(n_73), .ZN(n_0_151));
   OAI21_X1 i_0_282 (.A(n_0_153), .B1(n_0_199), .B2(n_0_274), .ZN(n_0_152));
   AOI21_X1 i_0_283 (.A(n_0_154), .B1(n_0_200), .B2(n_75), .ZN(n_0_153));
   NAND3_X1 i_0_284 (.A1(n_0_198), .A2(n_0_197), .A3(n_0_156), .ZN(n_0_154));
   NAND2_X1 i_0_285 (.A1(n_0_197), .A2(n_0_156), .ZN(n_0_155));
   OAI21_X1 i_0_286 (.A(n_0_200), .B1(n_0_157), .B2(n_78), .ZN(n_0_156));
   NAND2_X1 i_0_287 (.A1(n_0_160), .A2(n_0_273), .ZN(n_0_157));
   AOI21_X1 i_0_288 (.A(n_0_159), .B1(n_0_200), .B2(n_79), .ZN(n_0_158));
   NOR2_X1 i_0_289 (.A1(n_0_160), .A2(n_0_199), .ZN(n_0_159));
   NOR2_X1 i_0_290 (.A1(n_80), .A2(n_0_161), .ZN(n_0_160));
   INV_X1 i_0_291 (.A(n_0_162), .ZN(n_0_161));
   NAND3_X1 i_0_292 (.A1(n_0_174), .A2(n_0_169), .A3(n_0_163), .ZN(n_0_162));
   AOI21_X1 i_0_293 (.A(n_0_164), .B1(n_0_269), .B2(n_94), .ZN(n_0_163));
   NAND4_X1 i_0_294 (.A1(n_0_168), .A2(n_0_167), .A3(n_0_166), .A4(n_0_165), 
      .ZN(n_0_164));
   NOR4_X1 i_0_295 (.A1(n_87), .A2(n_90), .A3(n_91), .A4(n_93), .ZN(n_0_165));
   NOR3_X1 i_0_296 (.A1(n_88), .A2(n_89), .A3(n_92), .ZN(n_0_166));
   NOR4_X1 i_0_297 (.A1(n_83), .A2(n_84), .A3(n_85), .A4(n_86), .ZN(n_0_167));
   NOR2_X1 i_0_298 (.A1(n_81), .A2(n_82), .ZN(n_0_168));
   NAND4_X1 i_0_299 (.A1(n_0_173), .A2(n_0_172), .A3(n_0_171), .A4(n_0_170), 
      .ZN(n_0_169));
   NOR4_X1 i_0_300 (.A1(n_200), .A2(n_199), .A3(n_198), .A4(n_197), .ZN(n_0_170));
   NOR4_X1 i_0_301 (.A1(n_204), .A2(n_203), .A3(n_202), .A4(n_201), .ZN(n_0_171));
   NOR4_X1 i_0_302 (.A1(n_208), .A2(n_207), .A3(n_206), .A4(n_205), .ZN(n_0_172));
   NOR4_X1 i_0_303 (.A1(n_211), .A2(n_210), .A3(n_209), .A4(n_212), .ZN(n_0_173));
   OAI21_X1 i_0_304 (.A(n_0_175), .B1(n_0_177), .B2(n_0_176), .ZN(n_0_174));
   AOI22_X1 i_0_305 (.A1(n_211), .A2(n_0_69__1), .B1(n_0_74__1), .B2(n_212), 
      .ZN(n_0_175));
   OAI22_X1 i_0_306 (.A1(n_0_69__1), .A2(n_211), .B1(n_210), .B2(n_0_64__1), 
      .ZN(n_0_176));
   AOI221_X1 i_0_307 (.A(n_0_178), .B1(n_209), .B2(n_0_59__1), .C1(n_0_64__1), 
      .C2(n_210), .ZN(n_0_177));
   AOI21_X1 i_0_308 (.A(n_0_179), .B1(n_0_181), .B2(n_0_180), .ZN(n_0_178));
   OAI22_X1 i_0_309 (.A1(n_0_54__1), .A2(n_208), .B1(n_209), .B2(n_0_59__1), 
      .ZN(n_0_179));
   AOI22_X1 i_0_310 (.A1(n_0_54__1), .A2(n_208), .B1(n_207), .B2(n_0_49__1), 
      .ZN(n_0_180));
   OR2_X1 i_0_311 (.A1(n_0_183), .A2(n_0_182), .ZN(n_0_181));
   OAI22_X1 i_0_312 (.A1(n_207), .A2(n_0_49__1), .B1(n_0_44__1), .B2(n_206), 
      .ZN(n_0_182));
   AOI221_X1 i_0_313 (.A(n_0_184), .B1(n_205), .B2(n_0_39__1), .C1(n_0_44__1), 
      .C2(n_206), .ZN(n_0_183));
   AOI21_X1 i_0_314 (.A(n_0_185), .B1(n_0_187), .B2(n_0_186), .ZN(n_0_184));
   OAI22_X1 i_0_315 (.A1(n_0_34__1), .A2(n_204), .B1(n_205), .B2(n_0_39__1), 
      .ZN(n_0_185));
   AOI22_X1 i_0_316 (.A1(n_0_34__1), .A2(n_204), .B1(n_203), .B2(n_0_29__1), 
      .ZN(n_0_186));
   OR2_X1 i_0_317 (.A1(n_0_189), .A2(n_0_188), .ZN(n_0_187));
   OAI22_X1 i_0_318 (.A1(n_0_29__1), .A2(n_203), .B1(n_202), .B2(n_0_24__1), 
      .ZN(n_0_188));
   AOI21_X1 i_0_319 (.A(n_0_190), .B1(n_201), .B2(n_0_19__1), .ZN(n_0_189));
   OAI21_X1 i_0_320 (.A(n_0_191), .B1(n_0_193), .B2(n_0_192), .ZN(n_0_190));
   NAND2_X1 i_0_321 (.A1(n_202), .A2(n_0_24__1), .ZN(n_0_191));
   OAI22_X1 i_0_322 (.A1(n_0_19__1), .A2(n_201), .B1(n_200), .B2(n_0_14__1), 
      .ZN(n_0_192));
   AOI221_X1 i_0_323 (.A(n_0_194), .B1(n_199), .B2(n_0_9__1), .C1(n_0_14__1), 
      .C2(n_200), .ZN(n_0_193));
   AOI21_X1 i_0_324 (.A(n_0_195), .B1(n_0_196), .B2(n_109), .ZN(n_0_194));
   OAI22_X1 i_0_325 (.A1(n_0_9__1), .A2(n_199), .B1(n_198), .B2(n_0_4__1), 
      .ZN(n_0_195));
   AOI21_X1 i_0_326 (.A(n_197), .B1(n_198), .B2(n_0_4__1), .ZN(n_0_196));
   NAND2_X1 i_0_327 (.A1(n_77), .A2(n_0_200), .ZN(n_0_197));
   NAND2_X1 i_0_328 (.A1(n_76), .A2(n_0_200), .ZN(n_0_198));
   INV_X1 i_0_329 (.A(n_0_200), .ZN(n_0_199));
   AND2_X1 i_0_330 (.A1(n_65), .A2(n_0_205), .ZN(n_0_200));
   OAI21_X1 i_0_331 (.A(n_0_201), .B1(n_0_277), .B2(n_0), .ZN(n_193));
   NAND2_X1 i_0_332 (.A1(n_0_201), .A2(n_0), .ZN(QuotientVar[15]));
   NAND2_X1 i_0_333 (.A1(n_0_202), .A2(n_0_262), .ZN(n_0_201));
   XNOR2_X1 i_0_334 (.A(n_0_307), .B(Divisor[15]), .ZN(n_0_202));
   AOI21_X1 i_0_335 (.A(Reset), .B1(n_0_313), .B2(n_0_204), .ZN(n_194));
   NOR2_X1 i_0_336 (.A1(Reset), .A2(n_0_203), .ZN(n_195));
   NOR2_X1 i_0_337 (.A1(n_0_286), .A2(Start), .ZN(n_0_203));
   NAND2_X1 i_0_338 (.A1(n_0_205), .A2(n_0_286), .ZN(n_0_204));
   NOR3_X1 i_0_339 (.A1(n_0_206), .A2(n_32), .A3(n_31), .ZN(n_0_205));
   OR3_X1 i_0_340 (.A1(n_0_207), .A2(n_30), .A3(n_29), .ZN(n_0_206));
   INV_X1 i_0_341 (.A(n_0_208), .ZN(n_0_207));
   NOR3_X1 i_0_342 (.A1(n_0_218), .A2(n_0_213), .A3(n_0_209), .ZN(n_0_208));
   NAND3_X1 i_0_343 (.A1(n_0_212), .A2(n_0_211), .A3(n_0_210), .ZN(n_0_209));
   NOR2_X1 i_0_344 (.A1(n_11), .A2(n_12), .ZN(n_0_210));
   NOR2_X1 i_0_345 (.A1(n_9), .A2(n_10), .ZN(n_0_211));
   NOR4_X1 i_0_346 (.A1(n_13), .A2(n_14), .A3(n_15), .A4(n_16), .ZN(n_0_212));
   NAND4_X1 i_0_347 (.A1(n_0_217), .A2(n_0_216), .A3(n_0_215), .A4(n_0_214), 
      .ZN(n_0_213));
   NOR2_X1 i_0_348 (.A1(n_3), .A2(n_4), .ZN(n_0_214));
   NOR2_X1 i_0_349 (.A1(n_1), .A2(n_2), .ZN(n_0_215));
   NOR2_X1 i_0_350 (.A1(n_7), .A2(n_8), .ZN(n_0_216));
   NOR2_X1 i_0_351 (.A1(n_5), .A2(n_6), .ZN(n_0_217));
   NAND3_X1 i_0_352 (.A1(n_0_221), .A2(n_0_220), .A3(n_0_219), .ZN(n_0_218));
   NOR4_X1 i_0_353 (.A1(n_17), .A2(n_18), .A3(n_19), .A4(n_20), .ZN(n_0_219));
   NOR4_X1 i_0_354 (.A1(n_21), .A2(n_22), .A3(n_23), .A4(n_24), .ZN(n_0_220));
   NOR4_X1 i_0_355 (.A1(n_25), .A2(n_26), .A3(n_27), .A4(n_28), .ZN(n_0_221));
   OAI21_X1 i_0_356 (.A(n_0), .B1(n_0_222), .B2(n_0_313), .ZN(n_196));
   AND2_X1 i_0_357 (.A1(n_0_223), .A2(n_0_239), .ZN(n_0_222));
   OAI211_X1 i_0_358 (.A(n_0_245), .B(n_0_224), .C1(n_0_227), .C2(n_0_253), 
      .ZN(n_0_223));
   NOR2_X1 i_0_359 (.A1(n_0_20), .A2(n_0_1), .ZN(n_0_224));
   NOR3_X1 i_0_360 (.A1(n_0_226), .A2(Dividend[12]), .A3(Dividend[13]), .ZN(
      n_0_225));
   OAI21_X1 i_0_361 (.A(n_0_306), .B1(n_0_258), .B2(n_0_255), .ZN(n_0_226));
   NOR3_X1 i_0_362 (.A1(n_0_232), .A2(n_0_228), .A3(n_0_258), .ZN(n_0_227));
   AOI21_X1 i_0_363 (.A(Dividend[14]), .B1(n_0_229), .B2(n_0_256), .ZN(n_0_228));
   OAI211_X1 i_0_364 (.A(n_0_303), .B(n_0_302), .C1(n_0_230), .C2(n_0_255), 
      .ZN(n_0_229));
   AND3_X1 i_0_365 (.A1(n_0_299), .A2(n_0_298), .A3(n_0_231), .ZN(n_0_230));
   OAI211_X1 i_0_366 (.A(n_0_297), .B(n_0_296), .C1(Dividend[3]), .C2(
      Dividend[2]), .ZN(n_0_231));
   NAND2_X1 i_0_367 (.A1(n_0_306), .A2(n_0_233), .ZN(n_0_232));
   OAI21_X1 i_0_368 (.A(n_0_305), .B1(Dividend[12]), .B2(n_0_234), .ZN(n_0_233));
   AOI21_X1 i_0_369 (.A(Dividend[11]), .B1(n_0_302), .B2(n_0_235), .ZN(n_0_234));
   OAI21_X1 i_0_370 (.A(n_0_301), .B1(Dividend[8]), .B2(n_0_236), .ZN(n_0_235));
   AOI21_X1 i_0_371 (.A(Dividend[7]), .B1(n_0_298), .B2(n_0_237), .ZN(n_0_236));
   OAI21_X1 i_0_372 (.A(n_0_297), .B1(Dividend[4]), .B2(n_0_238), .ZN(n_0_237));
   AOI21_X1 i_0_373 (.A(Dividend[3]), .B1(n_0_294), .B2(Dividend[1]), .ZN(
      n_0_238));
   AOI21_X1 i_0_374 (.A(n_0_250), .B1(n_0_245), .B2(n_0_240), .ZN(n_0_239));
   AOI21_X1 i_0_375 (.A(n_0_241), .B1(Divisor[7]), .B2(Divisor[15]), .ZN(n_0_240));
   OR2_X1 i_0_376 (.A1(n_0_242), .A2(Divisor[6]), .ZN(n_0_241));
   OR3_X1 i_0_377 (.A1(n_0_243), .A2(Divisor[4]), .A3(Divisor[5]), .ZN(n_0_242));
   NAND3_X1 i_0_378 (.A1(n_0_244), .A2(n_0_287), .A3(n_0_288), .ZN(n_0_243));
   NOR2_X1 i_0_379 (.A1(Divisor[3]), .A2(Divisor[2]), .ZN(n_0_244));
   NOR3_X1 i_0_380 (.A1(n_0_247), .A2(n_0_246), .A3(Divisor[14]), .ZN(n_0_245));
   OR2_X1 i_0_381 (.A1(Divisor[13]), .A2(Divisor[12]), .ZN(n_0_246));
   NAND2_X1 i_0_382 (.A1(n_0_249), .A2(n_0_248), .ZN(n_0_247));
   NOR2_X1 i_0_383 (.A1(Divisor[9]), .A2(Divisor[8]), .ZN(n_0_248));
   NOR2_X1 i_0_384 (.A1(Divisor[11]), .A2(Divisor[10]), .ZN(n_0_249));
   NOR2_X1 i_0_385 (.A1(n_0_257), .A2(n_0_253), .ZN(n_0_250));
   NAND3_X1 i_0_386 (.A1(n_0_260), .A2(n_0_258), .A3(n_0_254), .ZN(n_0_251));
   NAND4_X1 i_0_387 (.A1(n_0_258), .A2(n_0_300), .A3(n_0_301), .A4(n_0_260), 
      .ZN(n_0_252));
   NAND3_X1 i_0_388 (.A1(n_0_254), .A2(n_0_306), .A3(n_0_256), .ZN(n_0_253));
   INV_X1 i_0_389 (.A(n_0_255), .ZN(n_0_254));
   NAND4_X1 i_0_390 (.A1(n_0_303), .A2(n_0_302), .A3(n_0_301), .A4(n_0_300), 
      .ZN(n_0_255));
   NOR2_X1 i_0_391 (.A1(Dividend[13]), .A2(Dividend[12]), .ZN(n_0_256));
   NAND2_X1 i_0_392 (.A1(n_0_260), .A2(n_0_258), .ZN(n_0_257));
   NOR4_X1 i_0_393 (.A1(Dividend[7]), .A2(Dividend[6]), .A3(Dividend[5]), 
      .A4(Dividend[4]), .ZN(n_0_258));
   NAND3_X1 i_0_394 (.A1(n_0_260), .A2(n_0_296), .A3(n_0_297), .ZN(n_0_259));
   INV_X1 i_0_395 (.A(n_0_261), .ZN(n_0_260));
   NAND4_X1 i_0_396 (.A1(n_0_295), .A2(n_0_294), .A3(n_0_293), .A4(n_0_292), 
      .ZN(n_0_261));
   AND2_X1 i_0_397 (.A1(Start), .A2(n_0), .ZN(n_0_262));
   AOI21_X1 i_0_398 (.A(n_0_263), .B1(n_126), .B2(n_0_278), .ZN(n_197));
   NOR2_X1 i_0_399 (.A1(n_125), .A2(n_126), .ZN(n_0_263));
   MUX2_X1 i_0_400 (.A(n_124), .B(addOut[1]), .S(n_126), .Z(n_198));
   MUX2_X1 i_0_401 (.A(n_123), .B(addOut[2]), .S(n_126), .Z(n_199));
   MUX2_X1 i_0_402 (.A(n_122), .B(addOut[3]), .S(n_126), .Z(n_200));
   AOI21_X1 i_0_403 (.A(n_0_264), .B1(n_126), .B2(n_0_279), .ZN(n_201));
   NOR2_X1 i_0_404 (.A1(n_121), .A2(n_126), .ZN(n_0_264));
   AOI21_X1 i_0_405 (.A(n_0_265), .B1(n_126), .B2(n_0_280), .ZN(n_202));
   NOR2_X1 i_0_406 (.A1(n_120), .A2(n_126), .ZN(n_0_265));
   MUX2_X1 i_0_407 (.A(n_119), .B(addOut[6]), .S(n_126), .Z(n_203));
   MUX2_X1 i_0_408 (.A(n_118), .B(addOut[7]), .S(n_126), .Z(n_204));
   AOI21_X1 i_0_409 (.A(n_0_266), .B1(n_126), .B2(n_0_281), .ZN(n_205));
   NOR2_X1 i_0_410 (.A1(n_117), .A2(n_126), .ZN(n_0_266));
   AOI21_X1 i_0_411 (.A(n_0_267), .B1(n_126), .B2(n_0_282), .ZN(n_206));
   NOR2_X1 i_0_412 (.A1(n_116), .A2(n_126), .ZN(n_0_267));
   MUX2_X1 i_0_413 (.A(n_115), .B(addOut[10]), .S(n_126), .Z(n_207));
   MUX2_X1 i_0_414 (.A(n_114), .B(addOut[11]), .S(n_126), .Z(n_208));
   AOI21_X1 i_0_415 (.A(n_0_268), .B1(n_126), .B2(n_0_283), .ZN(n_209));
   NOR2_X1 i_0_416 (.A1(n_113), .A2(n_126), .ZN(n_0_268));
   MUX2_X1 i_0_417 (.A(n_112), .B(addOut[13]), .S(n_126), .Z(n_210));
   MUX2_X1 i_0_418 (.A(n_111), .B(addOut[14]), .S(n_126), .Z(n_211));
   INV_X1 i_0_419 (.A(n_0_269), .ZN(n_212));
   OAI21_X1 i_0_420 (.A(n_0_270), .B1(n_126), .B2(n_110), .ZN(n_0_269));
   NAND2_X1 i_0_421 (.A1(n_0_284), .A2(n_126), .ZN(n_0_270));
   INV_X1 i_0_422 (.A(n_35), .ZN(n_0_271));
   INV_X1 i_0_423 (.A(n_37), .ZN(n_0_272));
   INV_X1 i_0_424 (.A(n_79), .ZN(n_0_273));
   INV_X1 i_0_425 (.A(n_74), .ZN(n_0_274));
   INV_X1 i_0_426 (.A(n_71), .ZN(n_0_275));
   INV_X1 i_0_427 (.A(n_68), .ZN(n_0_276));
   INV_X1 i_0_428 (.A(n_65), .ZN(n_0_277));
   INV_X1 i_0_429 (.A(addOut[0]), .ZN(n_0_278));
   INV_X1 i_0_430 (.A(addOut[4]), .ZN(n_0_279));
   INV_X1 i_0_431 (.A(addOut[5]), .ZN(n_0_280));
   INV_X1 i_0_432 (.A(addOut[8]), .ZN(n_0_281));
   INV_X1 i_0_433 (.A(addOut[9]), .ZN(n_0_282));
   INV_X1 i_0_434 (.A(addOut[12]), .ZN(n_0_283));
   INV_X1 i_0_435 (.A(addOut[15]), .ZN(n_0_284));
   INV_X1 i_0_436 (.A(Reset), .ZN(n_0_285));
   INV_X1 i_0_437 (.A(n_0), .ZN(n_0_286));
   INV_X1 i_0_438 (.A(Divisor[0]), .ZN(n_0_287));
   INV_X1 i_0_439 (.A(Divisor[1]), .ZN(n_0_288));
   INV_X1 i_0_440 (.A(Divisor[2]), .ZN(n_0_289));
   INV_X1 i_0_441 (.A(Divisor[10]), .ZN(n_0_290));
   INV_X1 i_0_442 (.A(Divisor[15]), .ZN(n_0_291));
   INV_X1 i_0_443 (.A(Dividend[0]), .ZN(n_0_292));
   INV_X1 i_0_444 (.A(Dividend[1]), .ZN(n_0_293));
   INV_X1 i_0_445 (.A(Dividend[2]), .ZN(n_0_294));
   INV_X1 i_0_446 (.A(Dividend[3]), .ZN(n_0_295));
   INV_X1 i_0_447 (.A(Dividend[4]), .ZN(n_0_296));
   INV_X1 i_0_448 (.A(Dividend[5]), .ZN(n_0_297));
   INV_X1 i_0_449 (.A(Dividend[6]), .ZN(n_0_298));
   INV_X1 i_0_450 (.A(Dividend[7]), .ZN(n_0_299));
   INV_X1 i_0_451 (.A(Dividend[8]), .ZN(n_0_300));
   INV_X1 i_0_452 (.A(Dividend[9]), .ZN(n_0_301));
   INV_X1 i_0_453 (.A(Dividend[10]), .ZN(n_0_302));
   INV_X1 i_0_454 (.A(Dividend[11]), .ZN(n_0_303));
   INV_X1 i_0_455 (.A(Dividend[12]), .ZN(n_0_304));
   INV_X1 i_0_456 (.A(Dividend[13]), .ZN(n_0_305));
   INV_X1 i_0_457 (.A(Dividend[14]), .ZN(n_0_306));
   INV_X1 i_0_458 (.A(Dividend[15]), .ZN(n_0_307));
   INV_X1 i_0_459 (.A(n_30), .ZN(n_0_308));
   INV_X1 i_0_460 (.A(n_109), .ZN(n_213));
   INV_X1 i_0_461 (.A(n_108), .ZN(n_0_4__1));
   INV_X1 i_0_462 (.A(n_107), .ZN(n_0_9__1));
   INV_X1 i_0_463 (.A(n_106), .ZN(n_0_14__1));
   INV_X1 i_0_464 (.A(n_105), .ZN(n_0_19__1));
   INV_X1 i_0_465 (.A(n_104), .ZN(n_0_24__1));
   INV_X1 i_0_466 (.A(n_103), .ZN(n_0_29__1));
   INV_X1 i_0_467 (.A(n_102), .ZN(n_0_34__1));
   INV_X1 i_0_468 (.A(n_101), .ZN(n_0_39__1));
   INV_X1 i_0_469 (.A(n_100), .ZN(n_0_44__1));
   INV_X1 i_0_470 (.A(n_99), .ZN(n_0_49__1));
   INV_X1 i_0_471 (.A(n_98), .ZN(n_0_54__1));
   INV_X1 i_0_472 (.A(n_97), .ZN(n_0_59__1));
   INV_X1 i_0_473 (.A(n_96), .ZN(n_0_64__1));
   INV_X1 i_0_474 (.A(n_95), .ZN(n_0_69__1));
   INV_X1 i_0_475 (.A(n_94), .ZN(n_0_74__1));
   INV_X1 i_0_476 (.A(n_92), .ZN(n_0_309));
   INV_X1 i_0_477 (.A(n_91), .ZN(n_0_310));
   INV_X1 i_0_478 (.A(n_89), .ZN(n_0_311));
   INV_X1 i_0_479 (.A(n_88), .ZN(n_0_312));
   INV_X1 i_0_480 (.A(n_0_262), .ZN(n_0_313));
endmodule

module Interpolation_Devision(Tk, Tz, Tn, CLK, reset, EN, Done, DivOut);
   input [15:0]Tk;
   input [15:0]Tz;
   input [15:0]Tn;
   input CLK;
   input reset;
   input EN;
   output Done;
   output [15:0]DivOut;

   wire [15:0]TkComp;
   wire [15:0]Tk_Tn;
   wire [15:0]Tz_Tn;
   wire Q2;
   wire Q1;
   wire DoneSignal;
   wire [15:0]Division_output;
   wire L1;
   wire [15:0]temp;
   wire n_16_3_0;
   wire n_16_3_1;
   wire n_16_3_2;

   TBUF_X1 i_0 (.A(Division_output[0]), .EN(n_0), .Z(DivOut[0]));
   TBUF_X1 i_1 (.A(Division_output[1]), .EN(n_0), .Z(DivOut[1]));
   TBUF_X1 i_2 (.A(Division_output[2]), .EN(n_0), .Z(DivOut[2]));
   TBUF_X1 i_3 (.A(Division_output[3]), .EN(n_0), .Z(DivOut[3]));
   TBUF_X1 i_4 (.A(Division_output[4]), .EN(n_0), .Z(DivOut[4]));
   TBUF_X1 i_5 (.A(Division_output[5]), .EN(n_0), .Z(DivOut[5]));
   TBUF_X1 i_6 (.A(Division_output[6]), .EN(n_0), .Z(DivOut[6]));
   TBUF_X1 i_7 (.A(Division_output[7]), .EN(n_0), .Z(DivOut[7]));
   TBUF_X1 i_8 (.A(Division_output[8]), .EN(n_0), .Z(DivOut[8]));
   TBUF_X1 i_9 (.A(Division_output[9]), .EN(n_0), .Z(DivOut[9]));
   TBUF_X1 i_10 (.A(Division_output[10]), .EN(n_0), .Z(DivOut[10]));
   TBUF_X1 i_11 (.A(Division_output[11]), .EN(n_0), .Z(DivOut[11]));
   TBUF_X1 i_12 (.A(Division_output[12]), .EN(n_0), .Z(DivOut[12]));
   TBUF_X1 i_13 (.A(Division_output[13]), .EN(n_0), .Z(DivOut[13]));
   TBUF_X1 i_14 (.A(Division_output[14]), .EN(n_0), .Z(DivOut[14]));
   TBUF_X1 i_15 (.A(Division_output[15]), .EN(n_0), .Z(DivOut[15]));
   Carry_Look_Ahead__0_467 add1 (.A(temp), .B(), .Cin(), .S({TkComp[15], 
      TkComp[14], TkComp[13], TkComp[12], TkComp[11], TkComp[10], TkComp[9], 
      TkComp[8], TkComp[7], TkComp[6], TkComp[5], TkComp[4], TkComp[3], 
      TkComp[2], TkComp[1], uc_0}));
   Carry_Look_Ahead__0_548 sub1 (.A(Tk), .B({TkComp[15], TkComp[14], TkComp[13], 
      TkComp[12], TkComp[11], TkComp[10], TkComp[9], TkComp[8], TkComp[7], 
      TkComp[6], TkComp[5], TkComp[4], TkComp[3], TkComp[2], TkComp[1], Tn[0]}), 
      .Cin(), .S(Tk_Tn));
   Carry_Look_Ahead__0_629 sub2 (.A(Tz), .B({TkComp[15], TkComp[14], TkComp[13], 
      TkComp[12], TkComp[11], TkComp[10], TkComp[9], TkComp[8], TkComp[7], 
      TkComp[6], TkComp[5], TkComp[4], TkComp[3], TkComp[2], TkComp[1], Tn[0]}), 
      .Cin(), .S(Tz_Tn));
   flipflop__0_835 F2 (.D(EN), .load(Q1), .Clk(CLK), .Q(Q2), .rst());
   flipflop F (.D(EN), .load(L1), .Clk(CLK), .Q(Q1), .rst(Q2));
   fixed_division D1 (.Dividend(Tk_Tn), .Divisor(Tz_Tn), .Reset(reset), .clk(), 
      .Start(Q1), .Quotient(Division_output), .ERR(), .Done(DoneSignal), 
      .OverFlow());
   INV_X1 i_16_0_0 (.A(reset), .ZN(L1));
   INV_X1 i_16_1_0 (.A(Tn[0]), .ZN(temp[0]));
   INV_X1 i_16_1_1 (.A(Tn[1]), .ZN(temp[1]));
   INV_X1 i_16_1_2 (.A(Tn[2]), .ZN(temp[2]));
   INV_X1 i_16_1_3 (.A(Tn[3]), .ZN(temp[3]));
   INV_X1 i_16_1_4 (.A(Tn[4]), .ZN(temp[4]));
   INV_X1 i_16_1_5 (.A(Tn[5]), .ZN(temp[5]));
   INV_X1 i_16_1_6 (.A(Tn[6]), .ZN(temp[6]));
   INV_X1 i_16_1_7 (.A(Tn[7]), .ZN(temp[7]));
   INV_X1 i_16_1_8 (.A(Tn[8]), .ZN(temp[8]));
   INV_X1 i_16_1_9 (.A(Tn[9]), .ZN(temp[9]));
   INV_X1 i_16_1_10 (.A(Tn[10]), .ZN(temp[10]));
   INV_X1 i_16_1_11 (.A(Tn[11]), .ZN(temp[11]));
   INV_X1 i_16_1_12 (.A(Tn[12]), .ZN(temp[12]));
   INV_X1 i_16_1_13 (.A(Tn[13]), .ZN(temp[13]));
   INV_X1 i_16_1_14 (.A(Tn[14]), .ZN(temp[14]));
   INV_X1 i_16_1_15 (.A(Tn[15]), .ZN(temp[15]));
   AND2_X1 i_16_2_0 (.A1(DoneSignal), .A2(EN), .ZN(Done));
   INV_X1 i_16_3_0 (.A(n_16_3_0), .ZN(n_0));
   NAND2_X1 i_16_3_1 (.A1(n_16_3_2), .A2(n_16_3_1), .ZN(n_16_3_0));
   INV_X1 i_16_3_2 (.A(DoneSignal), .ZN(n_16_3_1));
   INV_X1 i_16_3_3 (.A(EN), .ZN(n_16_3_2));
endmodule

module reg__0_811(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;

   DFF_X1 \Q_reg[15]  (.D(n_0), .CK(n_1), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_2), .CK(n_1), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_3), .CK(n_1), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_4), .CK(n_1), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_5), .CK(n_1), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_6), .CK(n_1), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_7), .CK(n_1), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_1), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_9), .CK(n_1), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_10), .CK(n_1), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_11), .CK(n_1), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_12), .CK(n_1), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_13), .CK(n_1), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_14), .CK(n_1), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_15), .CK(n_1), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_16), .CK(n_1), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(rst), .ZN(n_0_0));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(D[15]), .ZN(n_0));
   INV_X1 i_0_2 (.A(Clk), .ZN(n_1));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(D[14]), .ZN(n_2));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(D[13]), .ZN(n_3));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(D[12]), .ZN(n_4));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(D[11]), .ZN(n_5));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(D[10]), .ZN(n_6));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(D[9]), .ZN(n_7));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(D[8]), .ZN(n_8));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(D[7]), .ZN(n_9));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(D[6]), .ZN(n_10));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(D[5]), .ZN(n_11));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(D[4]), .ZN(n_12));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(D[3]), .ZN(n_13));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(D[2]), .ZN(n_14));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(D[1]), .ZN(n_15));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(D[0]), .ZN(n_16));
endmodule

module reg__0_831(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module \reg (D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_2_0;
   wire n_2_1;
   wire n_2_2;
   wire n_2_3;
   wire n_3_0;
   wire n_3_1;
   wire n_3_2;
   wire n_3_3;
   wire n_4_0;
   wire n_4_1;
   wire n_4_2;
   wire n_4_3;
   wire n_5_0;
   wire n_5_1;
   wire n_5_2;
   wire n_5_3;
   wire n_6_0;
   wire n_6_1;
   wire n_6_2;
   wire n_6_3;
   wire n_7_0;
   wire n_7_1;
   wire n_7_2;
   wire n_7_3;
   wire n_8_0;
   wire n_8_1;
   wire n_8_2;
   wire n_8_3;
   wire n_9_0;
   wire n_9_1;
   wire n_9_2;
   wire n_9_3;
   wire n_10_0;
   wire n_10_1;
   wire n_10_2;
   wire n_10_3;
   wire n_11_0;
   wire n_11_1;
   wire n_11_2;
   wire n_11_3;
   wire n_12_0;
   wire n_12_1;
   wire n_12_2;
   wire n_12_3;
   wire n_13_0;
   wire n_13_1;
   wire n_13_2;
   wire n_13_3;
   wire n_14_0;
   wire n_14_1;
   wire n_14_2;
   wire n_14_3;
   wire n_15_0;
   wire n_15_1;
   wire n_15_2;
   wire n_15_3;
   wire n_16_0;
   wire n_16_1;
   wire n_16_2;
   wire n_16_3;
   wire n_17_0;
   wire n_17_1;
   wire n_17_2;
   wire n_17_3;

   DFF_X1 \Q_reg[15]  (.D(n_10), .CK(n_1), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_11), .CK(n_1), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_12), .CK(n_1), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_13), .CK(n_1), .Q(Q[12]), .QN());
   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_0), .ZN(n_0));
   INV_X1 i_0_1 (.A(rst), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(load), .ZN(n_0_1));
   INV_X1 i_1_0 (.A(Clk), .ZN(n_1));
   INV_X1 i_2_0 (.A(n_0), .ZN(n_2_0));
   NAND2_X1 i_2_1 (.A1(n_2_0), .A2(Q[9]), .ZN(n_2_1));
   INV_X1 i_2_2 (.A(rst), .ZN(n_2_2));
   NAND2_X1 i_2_3 (.A1(D[9]), .A2(n_2_2), .ZN(n_2_3));
   OAI21_X1 i_2_4 (.A(n_2_1), .B1(n_2_3), .B2(n_2_0), .ZN(n_2));
   INV_X1 i_3_0 (.A(n_0), .ZN(n_3_0));
   NAND2_X1 i_3_1 (.A1(n_3_0), .A2(Q[6]), .ZN(n_3_1));
   INV_X1 i_3_2 (.A(rst), .ZN(n_3_2));
   NAND2_X1 i_3_3 (.A1(D[6]), .A2(n_3_2), .ZN(n_3_3));
   OAI21_X1 i_3_4 (.A(n_3_1), .B1(n_3_3), .B2(n_3_0), .ZN(n_3));
   INV_X1 i_4_0 (.A(n_0), .ZN(n_4_0));
   NAND2_X1 i_4_1 (.A1(n_4_0), .A2(Q[5]), .ZN(n_4_1));
   INV_X1 i_4_2 (.A(rst), .ZN(n_4_2));
   NAND2_X1 i_4_3 (.A1(D[5]), .A2(n_4_2), .ZN(n_4_3));
   OAI21_X1 i_4_4 (.A(n_4_1), .B1(n_4_3), .B2(n_4_0), .ZN(n_4));
   INV_X1 i_5_0 (.A(n_0), .ZN(n_5_0));
   NAND2_X1 i_5_1 (.A1(n_5_0), .A2(Q[4]), .ZN(n_5_1));
   INV_X1 i_5_2 (.A(rst), .ZN(n_5_2));
   NAND2_X1 i_5_3 (.A1(D[4]), .A2(n_5_2), .ZN(n_5_3));
   OAI21_X1 i_5_4 (.A(n_5_1), .B1(n_5_3), .B2(n_5_0), .ZN(n_5));
   INV_X1 i_6_0 (.A(n_0), .ZN(n_6_0));
   NAND2_X1 i_6_1 (.A1(n_6_0), .A2(Q[3]), .ZN(n_6_1));
   INV_X1 i_6_2 (.A(rst), .ZN(n_6_2));
   NAND2_X1 i_6_3 (.A1(D[3]), .A2(n_6_2), .ZN(n_6_3));
   OAI21_X1 i_6_4 (.A(n_6_1), .B1(n_6_3), .B2(n_6_0), .ZN(n_6));
   INV_X1 i_7_0 (.A(n_0), .ZN(n_7_0));
   NAND2_X1 i_7_1 (.A1(n_7_0), .A2(Q[2]), .ZN(n_7_1));
   INV_X1 i_7_2 (.A(rst), .ZN(n_7_2));
   NAND2_X1 i_7_3 (.A1(D[2]), .A2(n_7_2), .ZN(n_7_3));
   OAI21_X1 i_7_4 (.A(n_7_1), .B1(n_7_3), .B2(n_7_0), .ZN(n_7));
   INV_X1 i_8_0 (.A(n_0), .ZN(n_8_0));
   NAND2_X1 i_8_1 (.A1(n_8_0), .A2(Q[1]), .ZN(n_8_1));
   INV_X1 i_8_2 (.A(rst), .ZN(n_8_2));
   NAND2_X1 i_8_3 (.A1(D[1]), .A2(n_8_2), .ZN(n_8_3));
   OAI21_X1 i_8_4 (.A(n_8_1), .B1(n_8_3), .B2(n_8_0), .ZN(n_8));
   INV_X1 i_9_0 (.A(n_0), .ZN(n_9_0));
   NAND2_X1 i_9_1 (.A1(n_9_0), .A2(Q[0]), .ZN(n_9_1));
   INV_X1 i_9_2 (.A(rst), .ZN(n_9_2));
   NAND2_X1 i_9_3 (.A1(D[0]), .A2(n_9_2), .ZN(n_9_3));
   OAI21_X1 i_9_4 (.A(n_9_1), .B1(n_9_3), .B2(n_9_0), .ZN(n_9));
   NAND2_X1 i_10_0 (.A1(n_10_2), .A2(n_10_0), .ZN(n_10));
   NAND2_X1 i_10_1 (.A1(n_10_1), .A2(Q[15]), .ZN(n_10_0));
   INV_X1 i_10_2 (.A(n_0), .ZN(n_10_1));
   NAND3_X1 i_10_3 (.A1(D[15]), .A2(n_10_3), .A3(n_0), .ZN(n_10_2));
   INV_X1 i_10_4 (.A(rst), .ZN(n_10_3));
   NAND2_X1 i_11_0 (.A1(n_11_2), .A2(n_11_0), .ZN(n_11));
   NAND2_X1 i_11_1 (.A1(n_11_1), .A2(Q[14]), .ZN(n_11_0));
   INV_X1 i_11_2 (.A(n_0), .ZN(n_11_1));
   NAND3_X1 i_11_3 (.A1(D[14]), .A2(n_11_3), .A3(n_0), .ZN(n_11_2));
   INV_X1 i_11_4 (.A(rst), .ZN(n_11_3));
   NAND2_X1 i_12_0 (.A1(n_12_2), .A2(n_12_0), .ZN(n_12));
   NAND2_X1 i_12_1 (.A1(n_12_1), .A2(Q[13]), .ZN(n_12_0));
   INV_X1 i_12_2 (.A(n_0), .ZN(n_12_1));
   NAND3_X1 i_12_3 (.A1(D[13]), .A2(n_12_3), .A3(n_0), .ZN(n_12_2));
   INV_X1 i_12_4 (.A(rst), .ZN(n_12_3));
   NAND2_X1 i_13_0 (.A1(n_13_2), .A2(n_13_0), .ZN(n_13));
   NAND2_X1 i_13_1 (.A1(n_13_1), .A2(Q[12]), .ZN(n_13_0));
   INV_X1 i_13_2 (.A(n_0), .ZN(n_13_1));
   NAND3_X1 i_13_3 (.A1(D[12]), .A2(n_13_3), .A3(n_0), .ZN(n_13_2));
   INV_X1 i_13_4 (.A(rst), .ZN(n_13_3));
   NAND2_X1 i_14_0 (.A1(n_14_2), .A2(n_14_0), .ZN(n_14));
   NAND2_X1 i_14_1 (.A1(n_14_1), .A2(Q[11]), .ZN(n_14_0));
   INV_X1 i_14_2 (.A(n_0), .ZN(n_14_1));
   NAND3_X1 i_14_3 (.A1(D[11]), .A2(n_14_3), .A3(n_0), .ZN(n_14_2));
   INV_X1 i_14_4 (.A(rst), .ZN(n_14_3));
   NAND2_X1 i_15_0 (.A1(n_15_2), .A2(n_15_0), .ZN(n_15));
   NAND2_X1 i_15_1 (.A1(n_15_1), .A2(Q[10]), .ZN(n_15_0));
   INV_X1 i_15_2 (.A(n_0), .ZN(n_15_1));
   NAND3_X1 i_15_3 (.A1(D[10]), .A2(n_15_3), .A3(n_0), .ZN(n_15_2));
   INV_X1 i_15_4 (.A(rst), .ZN(n_15_3));
   NAND2_X1 i_16_0 (.A1(n_16_2), .A2(n_16_0), .ZN(n_16));
   NAND2_X1 i_16_1 (.A1(n_16_1), .A2(Q[8]), .ZN(n_16_0));
   INV_X1 i_16_2 (.A(n_0), .ZN(n_16_1));
   NAND3_X1 i_16_3 (.A1(D[8]), .A2(n_16_3), .A3(n_0), .ZN(n_16_2));
   INV_X1 i_16_4 (.A(rst), .ZN(n_16_3));
   NAND2_X1 i_17_0 (.A1(n_17_2), .A2(n_17_0), .ZN(n_17));
   NAND2_X1 i_17_1 (.A1(n_17_1), .A2(Q[7]), .ZN(n_17_0));
   INV_X1 i_17_2 (.A(n_0), .ZN(n_17_1));
   NAND3_X1 i_17_3 (.A1(D[7]), .A2(n_17_3), .A3(n_0), .ZN(n_17_2));
   INV_X1 i_17_4 (.A(rst), .ZN(n_17_3));
   DFF_X1 \Q_reg[11]  (.D(n_14), .CK(n_1), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_15), .CK(n_1), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_16), .CK(n_1), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_17), .CK(n_1), .Q(Q[7]), .QN());
   DFF_X2 \Q_reg[9]  (.D(n_2), .CK(n_1), .Q(Q[9]), .QN());
   DFF_X2 \Q_reg[5]  (.D(n_4), .CK(n_1), .Q(Q[5]), .QN());
   DFF_X2 \Q_reg[6]  (.D(n_3), .CK(n_1), .Q(Q[6]), .QN());
   DFF_X2 \Q_reg[3]  (.D(n_6), .CK(n_1), .Q(Q[3]), .QN());
   DFF_X2 \Q_reg[0]  (.D(n_9), .CK(n_1), .Q(Q[0]), .QN());
   DFF_X2 \Q_reg[4]  (.D(n_5), .CK(n_1), .Q(Q[4]), .QN());
   DFF_X2 \Q_reg[2]  (.D(n_7), .CK(n_1), .Q(Q[2]), .QN());
   DFF_X2 \Q_reg[1]  (.D(n_8), .CK(n_1), .Q(Q[1]), .QN());
endmodule

module Partial_Full_Adder__0_705(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_1_0;
   wire n_1_1;
   wire n_1_3;
   wire n_1_4;
   wire n_1_2;

   NAND2_X1 i_1_0 (.A1(A), .A2(Cin), .ZN(n_1_0));
   NAND2_X1 i_1_1 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_1));
   INV_X1 i_1_2 (.A(A), .ZN(n_1_3));
   INV_X1 i_1_3 (.A(Cin), .ZN(n_1_4));
   NAND2_X1 i_1_4 (.A1(n_1_0), .A2(n_1_1), .ZN(n_1_2));
   INV_X1 i_1_5 (.A(n_1_2), .ZN(S));
endmodule

module Partial_Full_Adder__0_701(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_697(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_693(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_689(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_685(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_681(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_677(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_673(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_669(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_665(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_661(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_657(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_653(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_649(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead__0_710(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire c15;
   wire c14;
   wire c13;
   wire c12;
   wire c11;
   wire c10;
   wire c9;
   wire c8;
   wire c7;
   wire c6;
   wire c5;
   wire c4;
   wire c3;
   wire c2;

   Partial_Full_Adder__0_705 PFA2 (.A(A[1]), .B(), .Cin(A[0]), .S(S[1]), .P(), 
      .G());
   Partial_Full_Adder__0_701 PFA3 (.A(A[2]), .B(), .Cin(c2), .S(S[2]), .P(), 
      .G());
   Partial_Full_Adder__0_697 PFA4 (.A(A[3]), .B(), .Cin(c3), .S(S[3]), .P(), 
      .G());
   Partial_Full_Adder__0_693 PFA5 (.A(A[4]), .B(), .Cin(c4), .S(S[4]), .P(), 
      .G());
   Partial_Full_Adder__0_689 PFA6 (.A(A[5]), .B(), .Cin(c5), .S(S[5]), .P(), 
      .G());
   Partial_Full_Adder__0_685 PFA7 (.A(A[6]), .B(), .Cin(c6), .S(S[6]), .P(), 
      .G());
   Partial_Full_Adder__0_681 PFA8 (.A(A[7]), .B(), .Cin(c7), .S(S[7]), .P(), 
      .G());
   Partial_Full_Adder__0_677 PFA9 (.A(A[8]), .B(), .Cin(c8), .S(S[8]), .P(), 
      .G());
   Partial_Full_Adder__0_673 PFA10 (.A(A[9]), .B(), .Cin(c9), .S(S[9]), .P(), 
      .G());
   Partial_Full_Adder__0_669 PFA11 (.A(A[10]), .B(), .Cin(c10), .S(S[10]), .P(), 
      .G());
   Partial_Full_Adder__0_665 PFA12 (.A(A[11]), .B(), .Cin(c11), .S(S[11]), .P(), 
      .G());
   Partial_Full_Adder__0_661 PFA13 (.A(A[12]), .B(), .Cin(c12), .S(S[12]), .P(), 
      .G());
   Partial_Full_Adder__0_657 PFA14 (.A(A[13]), .B(), .Cin(c13), .S(S[13]), .P(), 
      .G());
   Partial_Full_Adder__0_653 PFA15 (.A(A[14]), .B(), .Cin(c14), .S(S[14]), .P(), 
      .G());
   Partial_Full_Adder__0_649 PFA16 (.A(A[15]), .B(), .Cin(c15), .S(S[15]), .P(), 
      .G());
   AND2_X1 i_0_0 (.A1(A[14]), .A2(c14), .ZN(c15));
   AND2_X1 i_0_1 (.A1(A[13]), .A2(c13), .ZN(c14));
   AND2_X1 i_0_2 (.A1(A[12]), .A2(c12), .ZN(c13));
   AND2_X1 i_0_3 (.A1(A[11]), .A2(c11), .ZN(c12));
   AND2_X1 i_0_4 (.A1(A[10]), .A2(c10), .ZN(c11));
   AND2_X1 i_0_5 (.A1(A[9]), .A2(c9), .ZN(c10));
   AND2_X1 i_0_6 (.A1(A[8]), .A2(c8), .ZN(c9));
   AND2_X1 i_0_7 (.A1(A[7]), .A2(c7), .ZN(c8));
   AND2_X1 i_0_8 (.A1(A[6]), .A2(c6), .ZN(c7));
   AND2_X1 i_0_9 (.A1(A[5]), .A2(c5), .ZN(c6));
   AND2_X1 i_0_10 (.A1(A[4]), .A2(c4), .ZN(c5));
   AND2_X1 i_0_11 (.A1(A[3]), .A2(c3), .ZN(c4));
   AND2_X1 i_0_12 (.A1(A[2]), .A2(c2), .ZN(c3));
   AND2_X1 i_0_13 (.A1(A[0]), .A2(A[1]), .ZN(c2));
endmodule

module Partial_Full_Adder__0_790(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   NAND2_X1 i_0_0 (.A1(B), .A2(A), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(A), .ZN(n_0_2));
   INV_X1 i_0_3 (.A(B), .ZN(n_0_3));
   NAND2_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .ZN(n_0_4));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(S));
   AND2_X1 i_1_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_786(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_6;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_7;
   wire n_0_8;
   wire n_1_0;
   wire n_1_1;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
   INV_X1 i_0_0 (.A(Cin), .ZN(n_0_6));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(S));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(B), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_7), .A2(n_0_4), .ZN(n_0_2));
   NAND3_X1 i_0_5 (.A1(n_0_8), .A2(n_0_7), .A3(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(Cin), .A2(n_0_5), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(A), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_6), .A2(A), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(B), .ZN(n_0_8));
   INV_X1 i_1_0 (.A(B), .ZN(n_1_0));
   INV_X1 i_1_1 (.A(A), .ZN(n_1_1));
   OAI22_X1 i_1_2 (.A1(n_1_0), .A2(A), .B1(B), .B2(n_1_1), .ZN(P));
endmodule

module Partial_Full_Adder__0_782(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_778(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_774(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_770(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_766(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_762(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_758(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_754(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_750(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_746(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_742(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_738(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_734(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_730(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead__0_791(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire c1;
   wire c15;
   wire n_0_0;
   wire c14;
   wire n_0_1;
   wire c13;
   wire n_0_2;
   wire c12;
   wire n_0_3;
   wire c11;
   wire n_0_4;
   wire c10;
   wire n_0_5;
   wire c9;
   wire n_0_6;
   wire c8;
   wire n_0_7;
   wire c7;
   wire n_0_8;
   wire c6;
   wire n_0_9;
   wire c5;
   wire n_0_10;
   wire c4;
   wire n_0_11;
   wire c3;
   wire n_0_12;
   wire c2;
   wire n_0_13;

   Partial_Full_Adder__0_790 PFA1 (.A(A[0]), .B(B[0]), .Cin(), .S(S[0]), .P(), 
      .G(c1));
   Partial_Full_Adder__0_786 PFA2 (.A(A[1]), .B(B[1]), .Cin(c1), .S(S[1]), 
      .P(n_1), .G(n_0));
   Partial_Full_Adder__0_782 PFA3 (.A(A[2]), .B(B[2]), .Cin(c2), .S(S[2]), 
      .P(n_3), .G(n_2));
   Partial_Full_Adder__0_778 PFA4 (.A(A[3]), .B(B[3]), .Cin(c3), .S(S[3]), 
      .P(n_5), .G(n_4));
   Partial_Full_Adder__0_774 PFA5 (.A(A[4]), .B(B[4]), .Cin(c4), .S(S[4]), 
      .P(n_7), .G(n_6));
   Partial_Full_Adder__0_770 PFA6 (.A(A[5]), .B(B[5]), .Cin(c5), .S(S[5]), 
      .P(n_9), .G(n_8));
   Partial_Full_Adder__0_766 PFA7 (.A(A[6]), .B(B[6]), .Cin(c6), .S(S[6]), 
      .P(n_11), .G(n_10));
   Partial_Full_Adder__0_762 PFA8 (.A(A[7]), .B(B[7]), .Cin(c7), .S(S[7]), 
      .P(n_13), .G(n_12));
   Partial_Full_Adder__0_758 PFA9 (.A(A[8]), .B(B[8]), .Cin(c8), .S(S[8]), 
      .P(n_15), .G(n_14));
   Partial_Full_Adder__0_754 PFA10 (.A(A[9]), .B(B[9]), .Cin(c9), .S(S[9]), 
      .P(n_17), .G(n_16));
   Partial_Full_Adder__0_750 PFA11 (.A(A[10]), .B(B[10]), .Cin(c10), .S(S[10]), 
      .P(n_19), .G(n_18));
   Partial_Full_Adder__0_746 PFA12 (.A(A[11]), .B(B[11]), .Cin(c11), .S(S[11]), 
      .P(n_21), .G(n_20));
   Partial_Full_Adder__0_742 PFA13 (.A(A[12]), .B(B[12]), .Cin(c12), .S(S[12]), 
      .P(n_23), .G(n_22));
   Partial_Full_Adder__0_738 PFA14 (.A(A[13]), .B(B[13]), .Cin(c13), .S(S[13]), 
      .P(n_25), .G(n_24));
   Partial_Full_Adder__0_734 PFA15 (.A(A[14]), .B(B[14]), .Cin(c14), .S(S[14]), 
      .P(n_27), .G(n_26));
   Partial_Full_Adder__0_730 PFA16 (.A(A[15]), .B(B[15]), .Cin(c15), .S(S[15]), 
      .P(), .G());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(c15));
   AOI21_X1 i_0_1 (.A(n_26), .B1(n_27), .B2(c14), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(c14));
   AOI21_X1 i_0_3 (.A(n_24), .B1(n_25), .B2(c13), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(c13));
   AOI21_X1 i_0_5 (.A(n_22), .B1(n_23), .B2(c12), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(c12));
   AOI21_X1 i_0_7 (.A(n_20), .B1(n_21), .B2(c11), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(c11));
   AOI21_X1 i_0_9 (.A(n_18), .B1(n_19), .B2(c10), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(c10));
   AOI21_X1 i_0_11 (.A(n_16), .B1(n_17), .B2(c9), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(c9));
   AOI21_X1 i_0_13 (.A(n_14), .B1(n_15), .B2(c8), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(c8));
   AOI21_X1 i_0_15 (.A(n_12), .B1(n_13), .B2(c7), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(c7));
   AOI21_X1 i_0_17 (.A(n_10), .B1(n_11), .B2(c6), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(c6));
   AOI21_X1 i_0_19 (.A(n_8), .B1(n_9), .B2(c5), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(c5));
   AOI21_X1 i_0_21 (.A(n_6), .B1(n_7), .B2(c4), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(c4));
   AOI21_X1 i_0_23 (.A(n_4), .B1(n_5), .B2(c3), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(c3));
   AOI21_X1 i_0_25 (.A(n_2), .B1(n_3), .B2(c2), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(c2));
   AOI21_X1 i_0_27 (.A(n_0), .B1(c1), .B2(n_1), .ZN(n_0_13));
endmodule

module datapath__2_486(R, L, plus);
   input [32:0]R;
   input [32:0]L;
   output [32:0]plus;

   INV_X1 i_0 (.A(L[27]), .ZN(n_0));
   INV_X1 i_1 (.A(R[27]), .ZN(n_1));
   INV_X1 i_2 (.A(R[17]), .ZN(n_2));
   XNOR2_X1 i_3 (.A(L[17]), .B(n_2), .ZN(plus[17]));
   INV_X1 i_6 (.A(n_45), .ZN(n_4));
   OAI21_X1 i_7 (.A(n_100), .B1(n_12), .B2(n_4), .ZN(n_5));
   INV_X1 i_8 (.A(n_84), .ZN(n_6));
   NAND2_X1 i_9 (.A1(L[27]), .A2(R[27]), .ZN(n_7));
   NAND3_X1 i_11 (.A1(n_42), .A2(n_84), .A3(n_79), .ZN(n_9));
   NAND2_X1 i_12 (.A1(n_9), .A2(n_39), .ZN(n_10));
   NAND2_X1 i_10 (.A1(n_0), .A2(n_1), .ZN(n_11));
   NAND2_X1 i_14 (.A1(n_49), .A2(n_44), .ZN(n_12));
   AOI22_X1 i_13 (.A1(n_7), .A2(n_33), .B1(n_0), .B2(n_1), .ZN(n_14));
   OAI21_X1 i_16 (.A(n_39), .B1(n_105), .B2(n_34), .ZN(n_33));
   NAND2_X1 i_24 (.A1(L[28]), .A2(n_76), .ZN(n_16));
   NAND2_X1 i_26 (.A1(n_75), .A2(R[28]), .ZN(n_18));
   NAND2_X1 i_27 (.A1(L[28]), .A2(R[28]), .ZN(n_19));
   NAND2_X1 i_30 (.A1(n_75), .A2(n_76), .ZN(n_20));
   INV_X1 i_32 (.A(L[28]), .ZN(n_75));
   INV_X1 i_88 (.A(R[28]), .ZN(n_76));
   NAND2_X1 i_37 (.A1(n_11), .A2(n_78), .ZN(n_24));
   NAND2_X1 i_38 (.A1(n_7), .A2(n_10), .ZN(n_78));
   BUF_X1 i_4 (.A(n_55), .Z(n_51));
   BUF_X1 i_5 (.A(n_67), .Z(n_44));
   BUF_X1 i_15 (.A(n_102), .Z(n_45));
   INV_X1 i_39 (.A(n_42), .ZN(n_34));
   XOR2_X1 i_17 (.A(n_51), .B(n_3), .Z(plus[18]));
   OR2_X1 i_18 (.A1(n_13), .A2(n_54), .ZN(n_3));
   INV_X1 i_19 (.A(n_58), .ZN(n_13));
   NAND2_X1 i_21 (.A1(n_41), .A2(n_65), .ZN(n_31));
   XNOR2_X1 i_25 (.A(n_103), .B(n_57), .ZN(plus[21]));
   XNOR2_X1 i_22 (.A(n_21), .B(n_50), .ZN(plus[23]));
   NAND2_X1 i_23 (.A1(n_96), .A2(n_25), .ZN(n_21));
   XNOR2_X1 i_33 (.A(n_85), .B(n_22), .ZN(plus[24]));
   AOI21_X1 i_34 (.A(n_93), .B1(n_5), .B2(n_25), .ZN(n_22));
   XOR2_X1 i_35 (.A(n_92), .B(n_36), .Z(plus[25]));
   XNOR2_X1 i_36 (.A(n_29), .B(n_105), .ZN(plus[26]));
   NAND2_X1 i_20 (.A1(n_86), .A2(n_40), .ZN(plus[27]));
   NAND4_X1 i_28 (.A1(n_43), .A2(n_80), .A3(n_39), .A4(n_38), .ZN(n_40));
   INV_X1 i_55 (.A(R[27]), .ZN(n_15));
   NAND2_X1 i_29 (.A1(n_46), .A2(R[27]), .ZN(n_43));
   INV_X1 i_31 (.A(L[27]), .ZN(n_46));
   NAND2_X1 i_40 (.A1(n_96), .A2(n_50), .ZN(n_17));
   NAND2_X1 i_43 (.A1(n_62), .A2(n_49), .ZN(n_50));
   NOR2_X1 i_41 (.A1(L[18]), .A2(R[18]), .ZN(n_54));
   NAND2_X1 i_42 (.A1(L[17]), .A2(R[17]), .ZN(n_55));
   NAND2_X1 i_44 (.A1(L[18]), .A2(R[18]), .ZN(n_58));
   INV_X1 i_46 (.A(n_65), .ZN(n_37));
   NAND2_X1 i_47 (.A1(L[19]), .A2(R[19]), .ZN(n_65));
   OR2_X1 i_48 (.A1(L[19]), .A2(R[19]), .ZN(n_41));
   NAND2_X1 i_49 (.A1(L[23]), .A2(R[23]), .ZN(n_25));
   INV_X1 i_101 (.A(R[25]), .ZN(n_61));
   NAND2_X1 i_45 (.A1(n_53), .A2(n_100), .ZN(n_62));
   NAND2_X1 i_52 (.A1(n_102), .A2(n_67), .ZN(n_53));
   AOI21_X1 i_94 (.A(n_54), .B1(n_58), .B2(n_55), .ZN(n_73));
   XNOR2_X1 i_95 (.A(n_31), .B(n_73), .ZN(plus[19]));
   AOI21_X1 i_50 (.A(n_54), .B1(n_58), .B2(n_55), .ZN(n_60));
   NOR2_X1 i_53 (.A1(L[20]), .A2(R[20]), .ZN(n_52));
   NAND2_X1 i_71 (.A1(n_99), .A2(n_61), .ZN(n_26));
   NAND2_X1 i_51 (.A1(L[25]), .A2(R[25]), .ZN(n_89));
   INV_X1 i_107 (.A(n_61), .ZN(n_91));
   OAI21_X1 i_56 (.A(n_89), .B1(L[25]), .B2(n_91), .ZN(n_92));
   NOR2_X1 i_84 (.A1(L[23]), .A2(R[23]), .ZN(n_93));
   INV_X1 i_57 (.A(L[23]), .ZN(n_94));
   INV_X1 i_109 (.A(R[23]), .ZN(n_95));
   NAND2_X1 i_58 (.A1(n_94), .A2(n_95), .ZN(n_96));
   NAND3_X1 i_72 (.A1(n_20), .A2(n_19), .A3(n_24), .ZN(n_97));
   NAND3_X1 i_75 (.A1(n_18), .A2(n_16), .A3(n_14), .ZN(n_98));
   NAND2_X1 i_77 (.A1(n_97), .A2(n_98), .ZN(plus[28]));
   AOI21_X1 i_60 (.A(n_52), .B1(n_23), .B2(n_35), .ZN(n_57));
   AOI21_X1 i_69 (.A(n_52), .B1(n_23), .B2(n_35), .ZN(n_64));
   NAND2_X1 i_54 (.A1(L[27]), .A2(n_15), .ZN(n_80));
   INV_X1 i_81 (.A(L[25]), .ZN(n_99));
   XNOR2_X1 i_74 (.A(L[26]), .B(R[26]), .ZN(n_29));
   NAND2_X1 i_61 (.A1(L[20]), .A2(R[20]), .ZN(n_35));
   XNOR2_X1 i_59 (.A(L[20]), .B(R[20]), .ZN(n_66));
   OAI211_X1 i_65 (.A(n_42), .B(n_79), .C1(n_30), .C2(n_87), .ZN(n_38));
   OR2_X1 i_76 (.A1(L[26]), .A2(R[26]), .ZN(n_39));
   NAND2_X1 i_78 (.A1(L[26]), .A2(R[26]), .ZN(n_42));
   INV_X1 i_79 (.A(n_6), .ZN(n_30));
   INV_X1 i_80 (.A(n_26), .ZN(n_87));
   XNOR2_X1 i_82 (.A(L[27]), .B(n_15), .ZN(n_48));
   OAI21_X1 i_87 (.A(L[26]), .B1(n_26), .B2(R[26]), .ZN(n_56));
   NAND2_X1 i_90 (.A1(n_26), .A2(R[26]), .ZN(n_63));
   NAND2_X1 i_98 (.A1(n_56), .A2(n_63), .ZN(n_68));
   NAND2_X1 i_99 (.A1(L[26]), .A2(R[26]), .ZN(n_69));
   NAND2_X1 i_108 (.A1(n_47), .A2(n_27), .ZN(n_70));
   INV_X1 i_111 (.A(n_70), .ZN(n_77));
   NOR2_X1 i_102 (.A1(n_6), .A2(n_77), .ZN(n_81));
   NAND2_X1 i_104 (.A1(n_69), .A2(n_81), .ZN(n_82));
   NAND2_X1 i_106 (.A1(n_68), .A2(n_82), .ZN(n_83));
   NAND2_X1 i_112 (.A1(n_48), .A2(n_83), .ZN(n_86));
   INV_X1 i_100 (.A(n_101), .ZN(n_100));
   NOR2_X1 i_116 (.A1(L[22]), .A2(R[22]), .ZN(n_101));
   NAND2_X1 i_103 (.A1(L[21]), .A2(R[21]), .ZN(n_67));
   XNOR2_X1 i_66 (.A(L[21]), .B(R[21]), .ZN(n_103));
   OAI21_X1 i_70 (.A(n_64), .B1(L[21]), .B2(R[21]), .ZN(n_71));
   NAND2_X1 i_92 (.A1(n_71), .A2(n_67), .ZN(n_74));
   OAI21_X1 i_105 (.A(n_64), .B1(L[21]), .B2(R[21]), .ZN(n_102));
   OAI21_X1 i_62 (.A(n_41), .B1(n_60), .B2(n_37), .ZN(n_8));
   XOR2_X1 i_64 (.A(n_8), .B(n_66), .Z(plus[20]));
   OAI21_X1 i_73 (.A(n_41), .B1(n_60), .B2(n_37), .ZN(n_23));
   OR2_X1 i_67 (.A1(L[24]), .A2(R[24]), .ZN(n_27));
   NAND2_X1 i_68 (.A1(L[24]), .A2(R[24]), .ZN(n_28));
   XNOR2_X1 i_117 (.A(L[24]), .B(R[24]), .ZN(n_85));
   INV_X1 i_63 (.A(n_74), .ZN(n_90));
   XNOR2_X1 i_96 (.A(n_72), .B(n_90), .ZN(plus[22]));
   NAND3_X1 i_83 (.A1(n_28), .A2(n_25), .A3(n_17), .ZN(n_32));
   NAND2_X1 i_85 (.A1(n_27), .A2(n_32), .ZN(n_36));
   NAND3_X1 i_86 (.A1(n_28), .A2(n_25), .A3(n_17), .ZN(n_47));
   NAND2_X1 i_89 (.A1(L[22]), .A2(R[22]), .ZN(n_49));
   INV_X1 i_93 (.A(R[22]), .ZN(n_59));
   XNOR2_X1 i_97 (.A(L[22]), .B(n_59), .ZN(n_72));
   NAND3_X1 i_113 (.A1(n_27), .A2(n_26), .A3(n_47), .ZN(n_79));
   NAND2_X1 i_91 (.A1(L[25]), .A2(R[25]), .ZN(n_84));
   NAND3_X1 i_110 (.A1(n_26), .A2(n_47), .A3(n_27), .ZN(n_88));
   NAND2_X1 i_114 (.A1(L[25]), .A2(R[25]), .ZN(n_104));
   NAND2_X1 i_115 (.A1(n_88), .A2(n_104), .ZN(n_105));
endmodule

module datapath__2_495(R, L, plus);
   input [32:0]R;
   input [32:0]L;
   output [32:0]plus;

   INV_X1 i_0 (.A(n_0), .ZN(plus[17]));
   XNOR2_X1 i_1 (.A(L[17]), .B(R[17]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_33), .B(n_1), .Z(plus[18]));
   NAND2_X1 i_3 (.A1(n_2), .A2(n_34), .ZN(n_1));
   INV_X1 i_4 (.A(n_35), .ZN(n_2));
   XNOR2_X1 i_5 (.A(n_47), .B(n_3), .ZN(plus[19]));
   XNOR2_X1 i_10 (.A(n_66), .B(n_31), .ZN(plus[21]));
   XNOR2_X1 i_14 (.A(L[22]), .B(R[22]), .ZN(n_8));
   NAND2_X1 i_6 (.A1(n_53), .A2(n_44), .ZN(plus[25]));
   INV_X1 i_29 (.A(R[25]), .ZN(n_9));
   INV_X1 i_16 (.A(L[25]), .ZN(n_10));
   NAND3_X1 i_15 (.A1(n_16), .A2(n_15), .A3(n_12), .ZN(n_11));
   OAI21_X1 i_11 (.A(n_64), .B1(L[23]), .B2(R[23]), .ZN(n_12));
   AOI21_X1 i_38 (.A(n_35), .B1(n_34), .B2(n_33), .ZN(n_3));
   NAND2_X1 i_41 (.A1(L[17]), .A2(R[17]), .ZN(n_33));
   NAND2_X1 i_42 (.A1(L[18]), .A2(R[18]), .ZN(n_34));
   NOR2_X1 i_43 (.A1(L[18]), .A2(R[18]), .ZN(n_35));
   INV_X1 i_25 (.A(n_46), .ZN(n_6));
   NAND2_X1 i_12 (.A1(L[23]), .A2(R[23]), .ZN(n_15));
   NAND2_X1 i_13 (.A1(L[24]), .A2(R[24]), .ZN(n_16));
   INV_X1 i_17 (.A(L[24]), .ZN(n_17));
   INV_X1 i_56 (.A(R[24]), .ZN(n_21));
   NAND2_X1 i_7 (.A1(n_50), .A2(n_4), .ZN(plus[20]));
   NAND3_X1 i_8 (.A1(n_40), .A2(n_5), .A3(n_19), .ZN(n_4));
   NAND2_X1 i_9 (.A1(n_48), .A2(n_49), .ZN(n_5));
   INV_X1 i_40 (.A(L[20]), .ZN(n_48));
   INV_X1 i_48 (.A(R[20]), .ZN(n_49));
   OAI21_X1 i_45 (.A(n_58), .B1(n_51), .B2(n_20), .ZN(n_50));
   INV_X1 i_49 (.A(n_19), .ZN(n_51));
   NAND2_X1 i_24 (.A1(L[20]), .A2(R[20]), .ZN(n_19));
   NOR2_X1 i_57 (.A1(L[20]), .A2(R[20]), .ZN(n_20));
   NAND2_X1 i_18 (.A1(n_12), .A2(n_15), .ZN(n_22));
   XNOR2_X1 i_19 (.A(n_22), .B(n_29), .ZN(plus[24]));
   INV_X1 i_39 (.A(R[23]), .ZN(n_25));
   XNOR2_X1 i_32 (.A(L[23]), .B(n_25), .ZN(n_26));
   NAND2_X1 i_33 (.A1(n_26), .A2(n_24), .ZN(n_27));
   XNOR2_X1 i_50 (.A(n_61), .B(L[23]), .ZN(n_30));
   OAI21_X1 i_51 (.A(n_27), .B1(n_30), .B2(n_24), .ZN(plus[23]));
   AOI21_X1 i_26 (.A(n_20), .B1(n_40), .B2(n_19), .ZN(n_31));
   NAND2_X1 i_28 (.A1(n_11), .A2(n_32), .ZN(n_45));
   NAND2_X1 i_30 (.A1(n_57), .A2(n_45), .ZN(n_53));
   NAND2_X1 i_31 (.A1(n_11), .A2(n_32), .ZN(n_37));
   NAND2_X1 i_35 (.A1(n_10), .A2(R[25]), .ZN(n_56));
   NAND2_X1 i_37 (.A1(n_39), .A2(n_56), .ZN(n_57));
   NAND2_X1 i_20 (.A1(n_17), .A2(n_21), .ZN(n_23));
   NAND2_X1 i_21 (.A1(n_23), .A2(n_16), .ZN(n_29));
   NAND2_X1 i_22 (.A1(n_17), .A2(n_21), .ZN(n_32));
   OAI21_X1 i_46 (.A(n_7), .B1(n_6), .B2(n_3), .ZN(n_38));
   OR2_X1 i_65 (.A1(L[19]), .A2(R[19]), .ZN(n_7));
   NAND2_X1 i_66 (.A1(L[19]), .A2(R[19]), .ZN(n_46));
   XNOR2_X1 i_44 (.A(L[19]), .B(R[19]), .ZN(n_47));
   NOR2_X1 i_55 (.A1(L[22]), .A2(R[22]), .ZN(n_60));
   XNOR2_X1 i_62 (.A(n_60), .B(R[23]), .ZN(n_61));
   AOI21_X1 i_63 (.A(n_65), .B1(L[22]), .B2(R[22]), .ZN(n_24));
   NAND2_X1 i_47 (.A1(L[22]), .A2(R[22]), .ZN(n_28));
   NOR2_X1 i_53 (.A1(L[22]), .A2(R[22]), .ZN(n_63));
   OAI21_X1 i_23 (.A(n_28), .B1(n_36), .B2(n_63), .ZN(n_64));
   NAND2_X1 i_70 (.A1(L[25]), .A2(n_9), .ZN(n_39));
   NAND2_X1 i_71 (.A1(n_10), .A2(R[25]), .ZN(n_41));
   INV_X1 i_52 (.A(n_37), .ZN(n_42));
   NAND2_X1 i_73 (.A1(L[25]), .A2(n_9), .ZN(n_43));
   NAND3_X1 i_74 (.A1(n_41), .A2(n_42), .A3(n_43), .ZN(n_44));
   NAND2_X1 i_58 (.A1(n_19), .A2(n_38), .ZN(n_54));
   INV_X1 i_59 (.A(n_20), .ZN(n_55));
   NAND2_X1 i_64 (.A1(n_54), .A2(n_55), .ZN(n_13));
   XNOR2_X1 i_54 (.A(n_8), .B(n_65), .ZN(plus[22]));
   AOI21_X1 i_69 (.A(n_62), .B1(n_59), .B2(n_13), .ZN(n_65));
   NAND2_X1 i_67 (.A1(n_13), .A2(n_59), .ZN(n_14));
   INV_X1 i_72 (.A(n_62), .ZN(n_18));
   NAND2_X1 i_75 (.A1(n_14), .A2(n_18), .ZN(n_36));
   OAI21_X1 i_60 (.A(n_7), .B1(n_6), .B2(n_3), .ZN(n_40));
   OAI21_X1 i_61 (.A(n_7), .B1(n_6), .B2(n_3), .ZN(n_52));
   INV_X1 i_76 (.A(n_52), .ZN(n_58));
   NAND2_X1 i_27 (.A1(L[21]), .A2(R[21]), .ZN(n_59));
   NOR2_X1 i_34 (.A1(L[21]), .A2(R[21]), .ZN(n_62));
   XNOR2_X1 i_36 (.A(L[21]), .B(R[21]), .ZN(n_66));
endmodule

module datapath__2_498(R, L, plus);
   input [32:0]R;
   input [32:0]L;
   output [32:0]plus;

   INV_X1 i_0 (.A(n_0), .ZN(plus[17]));
   XNOR2_X1 i_1 (.A(L[17]), .B(R[17]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_9), .B(n_1), .Z(plus[18]));
   NAND2_X1 i_3 (.A1(n_61), .A2(n_10), .ZN(n_1));
   XNOR2_X1 i_5 (.A(n_3), .B(n_55), .ZN(plus[19]));
   NAND2_X1 i_6 (.A1(n_4), .A2(n_23), .ZN(n_3));
   INV_X1 i_7 (.A(n_24), .ZN(n_4));
   XNOR2_X1 i_8 (.A(n_5), .B(n_17), .ZN(plus[20]));
   NAND2_X1 i_9 (.A1(n_27), .A2(n_26), .ZN(n_5));
   XOR2_X1 i_10 (.A(n_8), .B(n_47), .Z(plus[21]));
   XNOR2_X1 i_13 (.A(n_38), .B(n_22), .ZN(plus[22]));
   NAND2_X1 i_4 (.A1(n_31), .A2(n_54), .ZN(n_6));
   INV_X1 i_19 (.A(R[22]), .ZN(n_7));
   OAI21_X1 i_11 (.A(n_27), .B1(n_25), .B2(n_17), .ZN(n_8));
   AOI21_X1 i_12 (.A(n_24), .B1(n_23), .B2(n_58), .ZN(n_17));
   NAND2_X1 i_26 (.A1(L[17]), .A2(R[17]), .ZN(n_9));
   NAND2_X1 i_24 (.A1(L[18]), .A2(R[18]), .ZN(n_10));
   NAND2_X1 i_15 (.A1(L[19]), .A2(R[19]), .ZN(n_23));
   NOR2_X1 i_16 (.A1(L[19]), .A2(R[19]), .ZN(n_24));
   INV_X1 i_14 (.A(n_26), .ZN(n_25));
   NAND2_X1 i_18 (.A1(L[20]), .A2(R[20]), .ZN(n_26));
   INV_X1 i_17 (.A(n_28), .ZN(n_27));
   NOR2_X1 i_21 (.A1(L[20]), .A2(R[20]), .ZN(n_28));
   NAND2_X1 i_20 (.A1(n_33), .A2(n_34), .ZN(n_32));
   INV_X1 i_22 (.A(L[24]), .ZN(n_33));
   INV_X1 i_40 (.A(R[24]), .ZN(n_34));
   NAND2_X1 i_23 (.A1(L[23]), .A2(R[23]), .ZN(n_11));
   NAND2_X1 i_25 (.A1(n_52), .A2(n_41), .ZN(plus[24]));
   NAND3_X1 i_27 (.A1(n_6), .A2(n_32), .A3(n_30), .ZN(n_41));
   NAND2_X1 i_28 (.A1(n_45), .A2(n_46), .ZN(n_29));
   INV_X1 i_29 (.A(L[24]), .ZN(n_45));
   INV_X1 i_54 (.A(R[24]), .ZN(n_46));
   NAND2_X1 i_31 (.A1(L[24]), .A2(R[24]), .ZN(n_30));
   NAND2_X1 i_42 (.A1(n_20), .A2(n_7), .ZN(n_36));
   NAND2_X1 i_57 (.A1(L[22]), .A2(R[22]), .ZN(n_37));
   NAND2_X1 i_58 (.A1(n_36), .A2(n_37), .ZN(n_38));
   NAND2_X1 i_32 (.A1(L[21]), .A2(R[21]), .ZN(n_16));
   NOR2_X1 i_33 (.A1(L[21]), .A2(R[21]), .ZN(n_18));
   XNOR2_X1 i_30 (.A(L[21]), .B(R[21]), .ZN(n_47));
   NAND2_X1 i_34 (.A1(n_48), .A2(n_49), .ZN(plus[23]));
   INV_X1 i_36 (.A(n_6), .ZN(n_50));
   NAND2_X1 i_37 (.A1(n_29), .A2(n_30), .ZN(n_51));
   NAND2_X1 i_38 (.A1(n_50), .A2(n_51), .ZN(n_52));
   OAI21_X1 i_39 (.A(n_19), .B1(n_14), .B2(n_22), .ZN(n_13));
   NAND2_X1 i_43 (.A1(n_11), .A2(n_53), .ZN(n_31));
   OAI21_X1 i_44 (.A(n_19), .B1(n_14), .B2(n_22), .ZN(n_53));
   OR2_X1 i_45 (.A1(L[23]), .A2(R[23]), .ZN(n_15));
   NAND3_X1 i_46 (.A1(n_15), .A2(n_13), .A3(n_11), .ZN(n_48));
   OR2_X1 i_47 (.A1(L[23]), .A2(R[23]), .ZN(n_54));
   NAND2_X1 i_48 (.A1(n_20), .A2(n_7), .ZN(n_19));
   INV_X1 i_49 (.A(L[22]), .ZN(n_20));
   AOI21_X1 i_50 (.A(n_18), .B1(n_16), .B2(n_8), .ZN(n_22));
   XNOR2_X1 i_51 (.A(L[23]), .B(R[23]), .ZN(n_35));
   INV_X1 i_35 (.A(n_7), .ZN(n_39));
   NOR2_X1 i_52 (.A1(L[22]), .A2(n_39), .ZN(n_40));
   AOI21_X1 i_41 (.A(n_18), .B1(n_8), .B2(n_16), .ZN(n_42));
   INV_X1 i_53 (.A(n_42), .ZN(n_43));
   AOI21_X1 i_55 (.A(n_40), .B1(n_2), .B2(n_43), .ZN(n_44));
   NAND2_X1 i_56 (.A1(n_35), .A2(n_44), .ZN(n_49));
   AOI21_X1 i_63 (.A(n_21), .B1(n_10), .B2(n_9), .ZN(n_55));
   INV_X1 i_64 (.A(n_21), .ZN(n_56));
   NAND2_X1 i_65 (.A1(n_10), .A2(n_9), .ZN(n_57));
   NAND2_X1 i_66 (.A1(n_56), .A2(n_57), .ZN(n_58));
   NAND2_X1 i_59 (.A1(L[22]), .A2(R[22]), .ZN(n_2));
   NAND2_X1 i_60 (.A1(L[22]), .A2(R[22]), .ZN(n_12));
   INV_X1 i_61 (.A(n_12), .ZN(n_14));
   NOR2_X1 i_62 (.A1(L[18]), .A2(R[18]), .ZN(n_21));
   INV_X1 i_67 (.A(L[18]), .ZN(n_59));
   INV_X1 i_68 (.A(R[18]), .ZN(n_60));
   NAND2_X1 i_69 (.A1(n_59), .A2(n_60), .ZN(n_61));
endmodule

module datapath__2_752(R, L, plus);
   input [32:0]R;
   input [32:0]L;
   output [32:0]plus;

   INV_X1 i_0 (.A(R[17]), .ZN(n_0));
   XNOR2_X1 i_1 (.A(L[17]), .B(n_0), .ZN(plus[17]));
   XNOR2_X1 i_5 (.A(n_3), .B(n_29), .ZN(plus[19]));
   XNOR2_X1 i_6 (.A(L[19]), .B(R[19]), .ZN(n_3));
   XNOR2_X1 i_7 (.A(n_4), .B(n_27), .ZN(plus[20]));
   NAND2_X1 i_8 (.A1(n_36), .A2(n_35), .ZN(n_4));
   XOR2_X1 i_9 (.A(n_26), .B(n_55), .Z(plus[21]));
   XNOR2_X1 i_10 (.A(n_53), .B(n_58), .ZN(plus[23]));
   NAND2_X1 i_11 (.A1(n_61), .A2(n_13), .ZN(plus[24]));
   NAND4_X1 i_15 (.A1(n_16), .A2(n_50), .A3(n_9), .A4(n_11), .ZN(n_13));
   INV_X1 i_23 (.A(R[24]), .ZN(n_6));
   NAND2_X1 i_16 (.A1(n_17), .A2(R[24]), .ZN(n_16));
   INV_X1 i_17 (.A(L[24]), .ZN(n_17));
   INV_X1 i_12 (.A(L[23]), .ZN(n_7));
   INV_X1 i_28 (.A(R[23]), .ZN(n_18));
   NAND2_X1 i_19 (.A1(n_19), .A2(n_14), .ZN(n_9));
   NAND2_X1 i_13 (.A1(n_26), .A2(n_8), .ZN(n_5));
   OAI21_X1 i_22 (.A(n_36), .B1(n_27), .B2(n_34), .ZN(n_26));
   NOR2_X1 i_24 (.A1(n_28), .A2(n_33), .ZN(n_27));
   AOI21_X1 i_25 (.A(n_29), .B1(L[19]), .B2(R[19]), .ZN(n_28));
   AOI21_X1 i_26 (.A(n_32), .B1(n_31), .B2(n_30), .ZN(n_29));
   NOR2_X1 i_29 (.A1(L[19]), .A2(R[19]), .ZN(n_33));
   INV_X1 i_31 (.A(n_35), .ZN(n_34));
   NAND2_X1 i_32 (.A1(L[20]), .A2(R[20]), .ZN(n_35));
   OR2_X1 i_35 (.A1(L[20]), .A2(R[20]), .ZN(n_36));
   NAND2_X1 i_36 (.A1(L[21]), .A2(R[21]), .ZN(n_8));
   NAND2_X1 i_14 (.A1(L[23]), .A2(R[23]), .ZN(n_19));
   NAND2_X1 i_2 (.A1(n_1), .A2(n_45), .ZN(plus[18]));
   OAI21_X1 i_3 (.A(n_44), .B1(n_2), .B2(n_32), .ZN(n_1));
   INV_X1 i_4 (.A(n_31), .ZN(n_2));
   NOR2_X1 i_37 (.A1(L[18]), .A2(R[18]), .ZN(n_32));
   INV_X1 i_39 (.A(n_30), .ZN(n_44));
   NAND3_X1 i_40 (.A1(n_46), .A2(n_30), .A3(n_31), .ZN(n_45));
   NAND2_X1 i_38 (.A1(L[18]), .A2(R[18]), .ZN(n_31));
   NAND2_X1 i_53 (.A1(n_47), .A2(n_48), .ZN(n_46));
   INV_X1 i_54 (.A(L[18]), .ZN(n_47));
   INV_X1 i_55 (.A(R[18]), .ZN(n_48));
   NAND2_X1 i_41 (.A1(L[17]), .A2(R[17]), .ZN(n_30));
   OAI21_X1 i_27 (.A(n_22), .B1(n_24), .B2(n_21), .ZN(n_14));
   INV_X1 i_57 (.A(n_40), .ZN(n_24));
   INV_X1 i_58 (.A(R[22]), .ZN(n_15));
   NAND2_X1 i_34 (.A1(L[22]), .A2(R[22]), .ZN(n_40));
   NAND2_X1 i_30 (.A1(L[24]), .A2(n_6), .ZN(n_50));
   NAND2_X1 i_33 (.A1(L[24]), .A2(n_6), .ZN(n_10));
   NAND2_X1 i_18 (.A1(n_7), .A2(n_18), .ZN(n_43));
   NAND2_X1 i_20 (.A1(n_43), .A2(n_19), .ZN(n_53));
   NAND2_X1 i_21 (.A1(n_7), .A2(n_18), .ZN(n_11));
   NAND2_X1 i_43 (.A1(n_5), .A2(n_20), .ZN(n_12));
   OR2_X1 i_62 (.A1(L[21]), .A2(R[21]), .ZN(n_49));
   NAND2_X1 i_63 (.A1(n_49), .A2(n_8), .ZN(n_55));
   NAND2_X1 i_45 (.A1(n_25), .A2(n_15), .ZN(n_22));
   INV_X1 i_48 (.A(L[22]), .ZN(n_25));
   INV_X1 i_51 (.A(R[22]), .ZN(n_38));
   NAND2_X1 i_42 (.A1(n_37), .A2(n_38), .ZN(n_39));
   OAI211_X1 i_50 (.A(L[22]), .B(n_39), .C1(n_5), .C2(R[22]), .ZN(n_42));
   INV_X1 i_64 (.A(n_15), .ZN(n_56));
   NAND3_X1 i_44 (.A1(n_5), .A2(n_20), .A3(n_56), .ZN(n_57));
   NAND2_X1 i_46 (.A1(n_42), .A2(n_57), .ZN(n_58));
   OR2_X1 i_52 (.A1(L[21]), .A2(R[21]), .ZN(n_20));
   NOR2_X1 i_59 (.A1(L[21]), .A2(R[21]), .ZN(n_37));
   INV_X1 i_47 (.A(n_12), .ZN(n_21));
   INV_X1 i_49 (.A(R[22]), .ZN(n_23));
   XNOR2_X1 i_56 (.A(L[22]), .B(n_23), .ZN(n_41));
   XNOR2_X1 i_67 (.A(n_41), .B(n_12), .ZN(plus[22]));
   INV_X1 i_60 (.A(L[24]), .ZN(n_51));
   INV_X1 i_61 (.A(n_6), .ZN(n_52));
   NAND2_X1 i_65 (.A1(n_51), .A2(n_52), .ZN(n_54));
   NAND2_X1 i_66 (.A1(n_10), .A2(n_54), .ZN(n_59));
   NAND2_X1 i_68 (.A1(n_9), .A2(n_11), .ZN(n_60));
   NAND2_X1 i_69 (.A1(n_59), .A2(n_60), .ZN(n_61));
endmodule

module booth_multiplier(m, r, result, overflow);
   input [15:0]m;
   input [15:0]r;
   output [15:0]result;
   output overflow;

   wire n_2_0;
   wire n_2_1;
   wire n_2_2;
   wire n_2_3;
   wire n_2_4;
   wire n_2_5;
   wire n_2_6;
   wire n_2_7;
   wire n_2_8;
   wire n_2_9;
   wire n_2_10;
   wire n_2_11;
   wire n_2_12;
   wire n_2_13;
   wire n_2_14;
   wire n_2_15;
   wire n_2_16;
   wire n_2_17;
   wire n_2_18;
   wire n_2_19;
   wire n_2_20;
   wire n_2_21;
   wire n_2_22;
   wire n_2_23;
   wire n_2_24;
   wire n_2_25;
   wire n_2_26;
   wire n_2_27;
   wire n_2_28;
   wire n_2_29;
   wire n_2_30;
   wire n_2_31;
   wire n_2_32;
   wire n_2_33;
   wire n_2_34;
   wire n_2_35;
   wire n_45_0;
   wire n_45_1;
   wire n_45_2;
   wire n_45_3;
   wire n_45_4;
   wire n_45_5;
   wire n_45_6;
   wire n_45_7;
   wire n_45_8;
   wire n_45_9;
   wire n_0_8;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_5;
   wire n_0_1;
   wire n_0_2;
   wire n_0_7;
   wire n_0_20;
   wire n_0_18;
   wire n_0_21;
   wire n_0_24;
   wire n_0_28;
   wire n_0_29;
   wire n_0_0;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_35;
   wire n_0_42;
   wire n_0_43;
   wire n_0_46;
   wire n_0_47;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_3;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_26;
   wire n_0_15;
   wire n_0_22;
   wire n_0_41;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_74;
   wire n_0_75;
   wire n_0_77;
   wire n_0_9;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_23;
   wire n_0_27;
   wire n_0_93;
   wire n_0_97;
   wire n_0_98;
   wire n_0_44;
   wire n_0_61;
   wire n_0_62;
   wire n_0_108;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_63;
   wire n_0_64;
   wire n_0_72;
   wire n_0_17;
   wire n_0_73;
   wire n_0_99;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_79;
   wire n_0_139;
   wire n_0_140;
   wire n_0_100;
   wire n_0_80;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_155;
   wire n_0_82;
   wire n_0_157;
   wire n_0_90;
   wire n_0_4;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_91;
   wire n_0_6;
   wire n_0_175;
   wire n_0_179;
   wire n_0_95;
   wire n_0_70;
   wire n_0_16;
   wire n_0_45;
   wire n_0_94;
   wire n_0_103;
   wire n_0_104;
   wire n_0_165;
   wire n_0_166;
   wire n_0_181;
   wire n_0_96;
   wire n_0_30;
   wire n_0_81;
   wire n_0_186;
   wire n_0_159;
   wire n_0_102;
   wire n_0_105;
   wire n_0_118;
   wire n_0_122;
   wire n_0_48;
   wire n_0_124;
   wire n_0_76;
   wire n_0_136;
   wire n_0_161;
   wire n_0_162;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_156;
   wire n_0_158;
   wire n_0_106;
   wire n_0_109;
   wire n_0_119;
   wire n_0_120;
   wire n_0_123;
   wire n_0_154;
   wire n_0_19;
   wire n_0_25;
   wire n_0_160;
   wire n_0_173;
   wire n_0_180;
   wire n_0_182;
   wire n_0_184;
   wire n_0_188;
   wire n_0_189;
   wire n_0_134;
   wire n_0_138;
   wire n_0_177;
   wire n_0_176;
   wire n_0_174;
   wire n_0_185;
   wire n_0_187;
   wire n_0_163;
   wire n_0_135;
   wire n_0_125;
   wire n_0_126;
   wire n_0_71;
   wire n_0_92;
   wire n_0_101;
   wire n_0_137;
   wire n_0_147;
   wire n_0_164;
   wire n_0_183;
   wire n_0_191;
   wire n_0_192;
   wire n_0_194;
   wire n_0_195;
   wire n_0_10;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_54;
   wire n_0_110;
   wire n_0_130;
   wire n_0_141;
   wire n_0_69;
   wire n_0_201;
   wire n_0_193;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_78;
   wire n_0_83;
   wire n_0_196;
   wire n_0_200;
   wire n_0_211;
   wire n_0_107;
   wire n_0_121;
   wire n_0_178;
   wire n_0_190;
   wire n_0_142;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_5_0;
   wire n_5_1;
   wire n_5_2;
   wire n_5_3;
   wire n_5_4;
   wire n_5_5;
   wire n_5_6;
   wire n_5_7;
   wire n_5_8;
   wire n_5_9;
   wire n_5_10;
   wire n_5_11;
   wire n_5_13;
   wire n_5_17;
   wire n_5_18;
   wire n_5_19;
   wire n_5_20;
   wire n_5_21;
   wire n_5_23;
   wire n_5_22;
   wire n_5_24;
   wire n_5_30;
   wire n_5_31;
   wire n_5_32;
   wire n_5_33;
   wire n_5_34;
   wire n_5_35;
   wire n_5_25;
   wire n_5_39;
   wire n_5_14;
   wire n_5_41;
   wire n_5_42;
   wire n_5_15;
   wire n_5_44;
   wire n_5_45;
   wire n_5_46;
   wire n_5_12;
   wire n_5_4591;
   wire n_5_4592;
   wire n_5_40;
   wire n_5_4593;
   wire n_5_16;
   wire n_5_47;
   wire n_5_4595;
   wire n_5_48;
   wire n_5_4596;
   wire n_5_27;
   wire n_5_4598;
   wire n_5_37;
   wire n_5_49;
   wire n_5_4601;
   wire n_5_50;
   wire n_5_51;
   wire n_5_52;
   wire n_5_53;
   wire n_5_54;
   wire n_5_55;
   wire n_5_56;
   wire n_5_57;
   wire n_5_58;
   wire n_5_59;
   wire n_5_67;
   wire n_5_68;
   wire n_5_69;
   wire n_5_61;
   wire n_5_62;
   wire n_5_63;
   wire n_5_64;
   wire n_5_65;
   wire n_5_66;
   wire n_5_70;
   wire n_5_71;
   wire n_5_72;
   wire n_5_73;
   wire n_5_74;
   wire n_5_75;
   wire n_5_76;
   wire n_5_77;
   wire n_5_78;
   wire n_5_80;
   wire n_5_84;
   wire n_5_85;
   wire n_5_26;
   wire n_5_36;
   wire n_5_83;
   wire n_5_91;
   wire n_5_92;
   wire n_5_93;
   wire n_5_97;
   wire n_5_98;
   wire n_5_101;
   wire n_5_86;
   wire n_5_103;
   wire n_5_104;
   wire n_5_105;
   wire n_5_28;
   wire n_5_107;
   wire n_5_108;
   wire n_5_109;
   wire n_5_110;
   wire n_5_111;
   wire n_5_112;
   wire n_5_113;
   wire n_5_29;
   wire n_5_114;
   wire n_5_115;
   wire n_5_116;
   wire n_5_118;
   wire n_5_119;
   wire n_5_120;
   wire n_5_121;
   wire n_5_124;
   wire n_5_43;
   wire n_5_128;
   wire n_5_129;
   wire n_5_60;
   wire n_5_79;
   wire n_5_133;
   wire n_5_134;
   wire n_5_81;
   wire n_5_82;
   wire n_5_137;
   wire n_5_138;
   wire n_5_139;
   wire n_5_140;
   wire n_5_141;
   wire n_5_142;
   wire n_5_87;
   wire n_5_145;
   wire n_5_88;
   wire n_5_147;
   wire n_5_148;
   wire n_5_149;
   wire n_5_150;
   wire n_5_151;
   wire n_5_152;
   wire n_5_153;
   wire n_5_154;
   wire n_5_155;
   wire n_5_89;
   wire n_5_4606;
   wire n_5_161;
   wire n_5_3855;
   wire n_5_4607;
   wire n_5_100;
   wire n_5_117;
   wire n_5_4611;
   wire n_5_4612;
   wire n_5_38;
   wire n_5_4614;
   wire n_5_164;
   wire n_5_165;
   wire n_5_166;
   wire n_5_167;
   wire n_5_168;
   wire n_5_169;
   wire n_5_170;
   wire n_5_171;
   wire n_5_437;
   wire n_5_172;
   wire n_5_173;
   wire n_5_122;
   wire n_5_90;
   wire n_5_94;
   wire n_5_178;
   wire n_5_179;
   wire n_5_450;
   wire n_5_96;
   wire n_5_468;
   wire n_5_125;
   wire n_5_186;
   wire n_5_187;
   wire n_5_190;
   wire n_5_191;
   wire n_5_193;
   wire n_5_194;
   wire n_5_195;
   wire n_5_126;
   wire n_5_99;
   wire n_5_102;
   wire n_5_198;
   wire n_5_106;
   wire n_5_200;
   wire n_5_202;
   wire n_5_123;
   wire n_5_205;
   wire n_5_206;
   wire n_5_207;
   wire n_5_208;
   wire n_5_127;
   wire n_5_131;
   wire n_5_143;
   wire n_5_212;
   wire n_5_213;
   wire n_5_214;
   wire n_5_130;
   wire n_5_144;
   wire n_5_146;
   wire n_5_180;
   wire n_5_4620;
   wire n_5_4621;
   wire n_5_4622;
   wire n_5_132;
   wire n_5_3863;
   wire n_5_136;
   wire n_5_220;
   wire n_5_222;
   wire n_5_223;
   wire n_5_224;
   wire n_5_95;
   wire n_5_188;
   wire n_5_3866;
   wire n_5_227;
   wire n_5_3867;
   wire n_5_228;
   wire n_5_3868;
   wire n_5_229;
   wire n_5_3869;
   wire n_5_230;
   wire n_5_231;
   wire n_5_177;
   wire n_5_157;
   wire n_5_158;
   wire n_5_159;
   wire n_5_160;
   wire n_5_3877;
   wire n_5_3879;
   wire n_5_233;
   wire n_5_3880;
   wire n_5_234;
   wire n_5_235;
   wire n_5_236;
   wire n_5_237;
   wire n_5_238;
   wire n_5_135;
   wire n_5_3881;
   wire n_5_3882;
   wire n_5_3883;
   wire n_5_241;
   wire n_5_162;
   wire n_5_163;
   wire n_5_3886;
   wire n_5_3887;
   wire n_5_244;
   wire n_5_245;
   wire n_5_246;
   wire n_5_247;
   wire n_5_3888;
   wire n_5_3889;
   wire n_5_248;
   wire n_5_175;
   wire n_5_176;
   wire n_5_253;
   wire n_5_254;
   wire n_5_255;
   wire n_5_491;
   wire n_5_492;
   wire n_5_189;
   wire n_5_257;
   wire n_5_511;
   wire n_5_258;
   wire n_5_259;
   wire n_5_499;
   wire n_5_260;
   wire n_5_262;
   wire n_5_3893;
   wire n_5_264;
   wire n_5_181;
   wire n_5_266;
   wire n_5_267;
   wire n_5_268;
   wire n_5_269;
   wire n_5_512;
   wire n_5_271;
   wire n_5_272;
   wire n_5_273;
   wire n_5_274;
   wire n_5_275;
   wire n_5_276;
   wire n_5_502;
   wire n_5_277;
   wire n_5_278;
   wire n_5_279;
   wire n_5_3898;
   wire n_5_280;
   wire n_5_281;
   wire n_5_282;
   wire n_5_283;
   wire n_5_284;
   wire n_5_182;
   wire n_5_286;
   wire n_5_287;
   wire n_5_288;
   wire n_5_289;
   wire n_5_290;
   wire n_5_232;
   wire n_5_292;
   wire n_5_270;
   wire n_5_295;
   wire n_5_4626;
   wire n_5_296;
   wire n_5_297;
   wire n_5_298;
   wire n_5_299;
   wire n_5_3903;
   wire n_5_300;
   wire n_5_301;
   wire n_5_302;
   wire n_5_303;
   wire n_5_304;
   wire n_5_305;
   wire n_5_306;
   wire n_5_307;
   wire n_5_3904;
   wire n_5_3905;
   wire n_5_517;
   wire n_5_3906;
   wire n_5_3907;
   wire n_5_520;
   wire n_5_4627;
   wire n_5_3910;
   wire n_5_183;
   wire n_5_184;
   wire n_5_185;
   wire n_5_192;
   wire n_5_196;
   wire n_5_3916;
   wire n_5_324;
   wire n_5_217;
   wire n_5_329;
   wire n_5_218;
   wire n_5_3918;
   wire n_5_197;
   wire n_5_335;
   wire n_5_221;
   wire n_5_3920;
   wire n_5_350;
   wire n_5_343;
   wire n_5_351;
   wire n_5_344;
   wire n_5_345;
   wire n_5_545;
   wire n_5_3921;
   wire n_5_4631;
   wire n_5_360;
   wire n_5_361;
   wire n_5_225;
   wire n_5_226;
   wire n_5_369;
   wire n_5_370;
   wire n_5_242;
   wire n_5_243;
   wire n_5_249;
   wire n_5_250;
   wire n_5_379;
   wire n_5_251;
   wire n_5_459;
   wire n_5_383;
   wire n_5_384;
   wire n_5_385;
   wire n_5_386;
   wire n_5_4632;
   wire n_5_252;
   wire n_5_390;
   wire n_5_399;
   wire n_5_400;
   wire n_5_401;
   wire n_5_402;
   wire n_5_403;
   wire n_5_404;
   wire n_5_405;
   wire n_5_406;
   wire n_5_407;
   wire n_5_408;
   wire n_5_409;
   wire n_5_411;
   wire n_5_412;
   wire n_5_414;
   wire n_5_4633;
   wire n_5_4634;
   wire n_5_422;
   wire n_5_549;
   wire n_5_3927;
   wire n_5_550;
   wire n_5_428;
   wire n_5_261;
   wire n_5_430;
   wire n_5_199;
   wire n_5_433;
   wire n_5_3928;
   wire n_5_475;
   wire n_5_263;
   wire n_5_441;
   wire n_5_442;
   wire n_5_156;
   wire n_5_174;
   wire n_5_239;
   wire n_5_446;
   wire n_5_447;
   wire n_5_448;
   wire n_5_449;
   wire n_5_503;
   wire n_5_454;
   wire n_5_457;
   wire n_5_458;
   wire n_5_463;
   wire n_5_466;
   wire n_5_467;
   wire n_5_518;
   wire n_5_469;
   wire n_5_470;
   wire n_5_471;
   wire n_5_472;
   wire n_5_473;
   wire n_5_474;
   wire n_5_522;
   wire n_5_3934;
   wire n_5_477;
   wire n_5_478;
   wire n_5_479;
   wire n_5_554;
   wire n_5_496;
   wire n_5_484;
   wire n_5_485;
   wire n_5_507;
   wire n_5_308;
   wire n_5_494;
   wire n_5_508;
   wire n_5_309;
   wire n_5_265;
   wire n_5_556;
   wire n_5_4635;
   wire n_5_557;
   wire n_5_311;
   wire n_5_312;
   wire n_5_558;
   wire n_5_559;
   wire n_5_313;
   wire n_5_314;
   wire n_5_315;
   wire n_5_201;
   wire n_5_317;
   wire n_5_561;
   wire n_5_562;
   wire n_5_563;
   wire n_5_564;
   wire n_5_318;
   wire n_5_3938;
   wire n_5_565;
   wire n_5_319;
   wire n_5_320;
   wire n_5_321;
   wire n_5_322;
   wire n_5_328;
   wire n_5_330;
   wire n_5_3939;
   wire n_5_331;
   wire n_5_332;
   wire n_5_3940;
   wire n_5_337;
   wire n_5_338;
   wire n_5_339;
   wire n_5_340;
   wire n_5_341;
   wire n_5_568;
   wire n_5_342;
   wire n_5_285;
   wire n_5_3941;
   wire n_5_3942;
   wire n_5_348;
   wire n_5_349;
   wire n_5_352;
   wire n_5_3943;
   wire n_5_310;
   wire n_5_356;
   wire n_5_357;
   wire n_5_358;
   wire n_5_3944;
   wire n_5_359;
   wire n_5_362;
   wire n_5_323;
   wire n_5_366;
   wire n_5_571;
   wire n_5_368;
   wire n_5_572;
   wire n_5_371;
   wire n_5_346;
   wire n_5_380;
   wire n_5_382;
   wire n_5_365;
   wire n_5_388;
   wire n_5_389;
   wire n_5_203;
   wire n_5_209;
   wire n_5_577;
   wire n_5_391;
   wire n_5_325;
   wire n_5_326;
   wire n_5_392;
   wire n_5_393;
   wire n_5_394;
   wire n_5_395;
   wire n_5_396;
   wire n_5_397;
   wire n_5_398;
   wire n_5_327;
   wire n_5_3948;
   wire n_5_580;
   wire n_5_413;
   wire n_5_415;
   wire n_5_416;
   wire n_5_3949;
   wire n_5_417;
   wire n_5_423;
   wire n_5_424;
   wire n_5_3950;
   wire n_5_425;
   wire n_5_3951;
   wire n_5_426;
   wire n_5_3952;
   wire n_5_3953;
   wire n_5_427;
   wire n_5_3954;
   wire n_5_431;
   wire n_5_434;
   wire n_5_435;
   wire n_5_333;
   wire n_5_3957;
   wire n_5_590;
   wire n_5_591;
   wire n_5_210;
   wire n_5_4636;
   wire n_5_594;
   wire n_5_4637;
   wire n_5_597;
   wire n_5_334;
   wire n_5_336;
   wire n_5_529;
   wire n_5_603;
   wire n_5_3963;
   wire n_5_3964;
   wire n_5_607;
   wire n_5_608;
   wire n_5_609;
   wire n_5_610;
   wire n_5_617;
   wire n_5_3965;
   wire n_5_627;
   wire n_5_628;
   wire n_5_629;
   wire n_5_630;
   wire n_5_631;
   wire n_5_632;
   wire n_5_633;
   wire n_5_634;
   wire n_5_211;
   wire n_5_636;
   wire n_5_347;
   wire n_5_642;
   wire n_5_353;
   wire n_5_651;
   wire n_5_655;
   wire n_5_656;
   wire n_5_657;
   wire n_5_658;
   wire n_5_659;
   wire n_5_660;
   wire n_5_661;
   wire n_5_662;
   wire n_5_663;
   wire n_5_664;
   wire n_5_3967;
   wire n_5_666;
   wire n_5_668;
   wire n_5_3968;
   wire n_5_670;
   wire n_5_671;
   wire n_5_3969;
   wire n_5_675;
   wire n_5_354;
   wire n_5_679;
   wire n_5_682;
   wire n_5_683;
   wire n_5_355;
   wire n_5_685;
   wire n_5_686;
   wire n_5_687;
   wire n_5_688;
   wire n_5_3970;
   wire n_5_690;
   wire n_5_693;
   wire n_5_694;
   wire n_5_3971;
   wire n_5_696;
   wire n_5_4639;
   wire n_5_4640;
   wire n_5_3972;
   wire n_5_3973;
   wire n_5_710;
   wire n_5_363;
   wire n_5_592;
   wire n_5_712;
   wire n_5_713;
   wire n_5_3975;
   wire n_5_3976;
   wire n_5_444;
   wire n_5_3977;
   wire n_5_445;
   wire n_5_3979;
   wire n_5_4642;
   wire n_5_451;
   wire n_5_364;
   wire n_5_453;
   wire n_5_367;
   wire n_5_372;
   wire n_5_373;
   wire n_5_480;
   wire n_5_4644;
   wire n_5_481;
   wire n_5_482;
   wire n_5_483;
   wire n_5_3987;
   wire n_5_487;
   wire n_5_4645;
   wire n_5_488;
   wire n_5_489;
   wire n_5_490;
   wire n_5_3989;
   wire n_5_493;
   wire n_5_495;
   wire n_5_374;
   wire n_5_500;
   wire n_5_3990;
   wire n_5_501;
   wire n_5_504;
   wire n_5_505;
   wire n_5_3991;
   wire n_5_506;
   wire n_5_620;
   wire n_5_723;
   wire n_5_509;
   wire n_5_3993;
   wire n_5_510;
   wire n_5_513;
   wire n_5_4646;
   wire n_5_514;
   wire n_5_4647;
   wire n_5_375;
   wire n_5_516;
   wire n_5_3994;
   wire n_5_519;
   wire n_5_521;
   wire n_5_523;
   wire n_5_527;
   wire n_5_3996;
   wire n_5_4648;
   wire n_5_530;
   wire n_5_376;
   wire n_5_533;
   wire n_5_534;
   wire n_5_377;
   wire n_5_535;
   wire n_5_537;
   wire n_5_3998;
   wire n_5_538;
   wire n_5_540;
   wire n_5_541;
   wire n_5_542;
   wire n_5_543;
   wire n_5_544;
   wire n_5_547;
   wire n_5_3999;
   wire n_5_548;
   wire n_5_551;
   wire n_5_552;
   wire n_5_553;
   wire n_5_555;
   wire n_5_4001;
   wire n_5_4002;
   wire n_5_4003;
   wire n_5_560;
   wire n_5_566;
   wire n_5_567;
   wire n_5_569;
   wire n_5_4649;
   wire n_5_381;
   wire n_5_570;
   wire n_5_573;
   wire n_5_724;
   wire n_5_4005;
   wire n_5_4006;
   wire n_5_4007;
   wire n_5_574;
   wire n_5_575;
   wire n_5_410;
   wire n_5_418;
   wire n_5_419;
   wire n_5_582;
   wire n_5_583;
   wire n_5_4010;
   wire n_5_4011;
   wire n_5_4012;
   wire n_5_4013;
   wire n_5_420;
   wire n_5_378;
   wire n_5_4015;
   wire n_5_584;
   wire n_5_585;
   wire n_5_586;
   wire n_5_587;
   wire n_5_588;
   wire n_5_589;
   wire n_5_593;
   wire n_5_3332;
   wire n_5_595;
   wire n_5_596;
   wire n_5_598;
   wire n_5_599;
   wire n_5_3333;
   wire n_5_600;
   wire n_5_4653;
   wire n_5_601;
   wire n_5_604;
   wire n_5_605;
   wire n_5_606;
   wire n_5_611;
   wire n_5_612;
   wire n_5_4016;
   wire n_5_613;
   wire n_5_293;
   wire n_5_614;
   wire n_5_615;
   wire n_5_618;
   wire n_5_621;
   wire n_5_436;
   wire n_5_623;
   wire n_5_4017;
   wire n_5_3335;
   wire n_5_1006;
   wire n_5_624;
   wire n_5_635;
   wire n_5_637;
   wire n_5_638;
   wire n_5_639;
   wire n_5_640;
   wire n_5_4019;
   wire n_5_641;
   wire n_5_3338;
   wire n_5_4020;
   wire n_5_643;
   wire n_5_644;
   wire n_5_645;
   wire n_5_648;
   wire n_5_652;
   wire n_5_653;
   wire n_5_654;
   wire n_5_665;
   wire n_5_667;
   wire n_5_669;
   wire n_5_672;
   wire n_5_673;
   wire n_5_4021;
   wire n_5_674;
   wire n_5_676;
   wire n_5_677;
   wire n_5_680;
   wire n_5_681;
   wire n_5_3124;
   wire n_5_689;
   wire n_5_4022;
   wire n_5_691;
   wire n_5_695;
   wire n_5_697;
   wire n_5_698;
   wire n_5_699;
   wire n_5_703;
   wire n_5_3339;
   wire n_5_704;
   wire n_5_705;
   wire n_5_706;
   wire n_5_707;
   wire n_5_708;
   wire n_5_709;
   wire n_5_714;
   wire n_5_715;
   wire n_5_4023;
   wire n_5_4024;
   wire n_5_438;
   wire n_5_717;
   wire n_5_718;
   wire n_5_719;
   wire n_5_720;
   wire n_5_721;
   wire n_5_722;
   wire n_5_725;
   wire n_5_726;
   wire n_5_727;
   wire n_5_439;
   wire n_5_729;
   wire n_5_3126;
   wire n_5_730;
   wire n_5_731;
   wire n_5_732;
   wire n_5_3340;
   wire n_5_733;
   wire n_5_4025;
   wire n_5_734;
   wire n_5_735;
   wire n_5_736;
   wire n_5_737;
   wire n_5_3128;
   wire n_5_738;
   wire n_5_440;
   wire n_5_3129;
   wire n_5_740;
   wire n_5_741;
   wire n_5_742;
   wire n_5_743;
   wire n_5_744;
   wire n_5_4026;
   wire n_5_745;
   wire n_5_4027;
   wire n_5_4028;
   wire n_5_746;
   wire n_5_747;
   wire n_5_748;
   wire n_5_750;
   wire n_5_751;
   wire n_5_752;
   wire n_5_753;
   wire n_5_4029;
   wire n_5_754;
   wire n_5_755;
   wire n_5_756;
   wire n_5_757;
   wire n_5_758;
   wire n_5_759;
   wire n_5_760;
   wire n_5_761;
   wire n_5_762;
   wire n_5_763;
   wire n_5_764;
   wire n_5_765;
   wire n_5_766;
   wire n_5_767;
   wire n_5_768;
   wire n_5_769;
   wire n_5_770;
   wire n_5_771;
   wire n_5_772;
   wire n_5_3341;
   wire n_5_773;
   wire n_5_4030;
   wire n_5_4031;
   wire n_5_774;
   wire n_5_775;
   wire n_5_776;
   wire n_5_777;
   wire n_5_778;
   wire n_5_779;
   wire n_5_780;
   wire n_5_781;
   wire n_5_782;
   wire n_5_783;
   wire n_5_784;
   wire n_5_785;
   wire n_5_786;
   wire n_5_787;
   wire n_5_788;
   wire n_5_4032;
   wire n_5_789;
   wire n_5_790;
   wire n_5_3131;
   wire n_5_791;
   wire n_5_792;
   wire n_5_793;
   wire n_5_4033;
   wire n_5_794;
   wire n_5_795;
   wire n_5_796;
   wire n_5_797;
   wire n_5_798;
   wire n_5_799;
   wire n_5_800;
   wire n_5_801;
   wire n_5_802;
   wire n_5_803;
   wire n_5_804;
   wire n_5_805;
   wire n_5_806;
   wire n_5_807;
   wire n_5_808;
   wire n_5_809;
   wire n_5_4034;
   wire n_5_810;
   wire n_5_811;
   wire n_5_812;
   wire n_5_813;
   wire n_5_814;
   wire n_5_3343;
   wire n_5_815;
   wire n_5_816;
   wire n_5_817;
   wire n_5_818;
   wire n_5_819;
   wire n_5_820;
   wire n_5_452;
   wire n_5_822;
   wire n_5_3345;
   wire n_5_823;
   wire n_5_824;
   wire n_5_825;
   wire n_5_826;
   wire n_5_827;
   wire n_5_828;
   wire n_5_829;
   wire n_5_830;
   wire n_5_831;
   wire n_5_832;
   wire n_5_833;
   wire n_5_834;
   wire n_5_835;
   wire n_5_836;
   wire n_5_837;
   wire n_5_4035;
   wire n_5_838;
   wire n_5_839;
   wire n_5_840;
   wire n_5_841;
   wire n_5_4036;
   wire n_5_387;
   wire n_5_844;
   wire n_5_845;
   wire n_5_846;
   wire n_5_847;
   wire n_5_848;
   wire n_5_849;
   wire n_5_4038;
   wire n_5_4039;
   wire n_5_850;
   wire n_5_851;
   wire n_5_852;
   wire n_5_853;
   wire n_5_854;
   wire n_5_3136;
   wire n_5_855;
   wire n_5_856;
   wire n_5_857;
   wire n_5_3347;
   wire n_5_858;
   wire n_5_4041;
   wire n_5_859;
   wire n_5_860;
   wire n_5_4655;
   wire n_5_4042;
   wire n_5_861;
   wire n_5_862;
   wire n_5_863;
   wire n_5_864;
   wire n_5_865;
   wire n_5_4043;
   wire n_5_866;
   wire n_5_867;
   wire n_5_868;
   wire n_5_4044;
   wire n_5_869;
   wire n_5_870;
   wire n_5_871;
   wire n_5_872;
   wire n_5_3682;
   wire n_5_421;
   wire n_5_874;
   wire n_5_875;
   wire n_5_602;
   wire n_5_4045;
   wire n_5_877;
   wire n_5_842;
   wire n_5_879;
   wire n_5_3736;
   wire n_5_3808;
   wire n_5_880;
   wire n_5_881;
   wire n_5_882;
   wire n_5_883;
   wire n_5_884;
   wire n_5_885;
   wire n_5_886;
   wire n_5_887;
   wire n_5_888;
   wire n_5_889;
   wire n_5_890;
   wire n_5_891;
   wire n_5_892;
   wire n_5_893;
   wire n_5_894;
   wire n_5_895;
   wire n_5_896;
   wire n_5_897;
   wire n_5_898;
   wire n_5_899;
   wire n_5_900;
   wire n_5_901;
   wire n_5_902;
   wire n_5_903;
   wire n_5_3350;
   wire n_5_904;
   wire n_5_4048;
   wire n_5_4049;
   wire n_5_4050;
   wire n_5_905;
   wire n_5_3138;
   wire n_5_906;
   wire n_5_3139;
   wire n_5_4051;
   wire n_5_907;
   wire n_5_4052;
   wire n_5_4053;
   wire n_5_908;
   wire n_5_909;
   wire n_5_910;
   wire n_5_3352;
   wire n_5_911;
   wire n_5_455;
   wire n_5_912;
   wire n_5_913;
   wire n_5_914;
   wire n_5_915;
   wire n_5_916;
   wire n_5_917;
   wire n_5_918;
   wire n_5_919;
   wire n_5_920;
   wire n_5_921;
   wire n_5_922;
   wire n_5_4056;
   wire n_5_923;
   wire n_5_924;
   wire n_5_925;
   wire n_5_926;
   wire n_5_927;
   wire n_5_928;
   wire n_5_929;
   wire n_5_930;
   wire n_5_3141;
   wire n_5_931;
   wire n_5_932;
   wire n_5_933;
   wire n_5_1806;
   wire n_5_934;
   wire n_5_935;
   wire n_5_936;
   wire n_5_937;
   wire n_5_938;
   wire n_5_1817;
   wire n_5_1819;
   wire n_5_939;
   wire n_5_1820;
   wire n_5_940;
   wire n_5_3142;
   wire n_5_3143;
   wire n_5_941;
   wire n_5_942;
   wire n_5_943;
   wire n_5_3355;
   wire n_5_944;
   wire n_5_945;
   wire n_5_3356;
   wire n_5_3357;
   wire n_5_4057;
   wire n_5_3147;
   wire n_5_3148;
   wire n_5_946;
   wire n_5_947;
   wire n_5_3149;
   wire n_5_948;
   wire n_5_949;
   wire n_5_950;
   wire n_5_951;
   wire n_5_952;
   wire n_5_953;
   wire n_5_954;
   wire n_5_955;
   wire n_5_956;
   wire n_5_1826;
   wire n_5_1828;
   wire n_5_957;
   wire n_5_958;
   wire n_5_959;
   wire n_5_960;
   wire n_5_961;
   wire n_5_962;
   wire n_5_963;
   wire n_5_964;
   wire n_5_965;
   wire n_5_966;
   wire n_5_967;
   wire n_5_968;
   wire n_5_969;
   wire n_5_970;
   wire n_5_971;
   wire n_5_972;
   wire n_5_1844;
   wire n_5_973;
   wire n_5_974;
   wire n_5_975;
   wire n_5_976;
   wire n_5_1850;
   wire n_5_1863;
   wire n_5_977;
   wire n_5_978;
   wire n_5_979;
   wire n_5_980;
   wire n_5_981;
   wire n_5_982;
   wire n_5_983;
   wire n_5_984;
   wire n_5_985;
   wire n_5_986;
   wire n_5_987;
   wire n_5_988;
   wire n_5_3151;
   wire n_5_989;
   wire n_5_990;
   wire n_5_3152;
   wire n_5_991;
   wire n_5_992;
   wire n_5_993;
   wire n_5_994;
   wire n_5_995;
   wire n_5_3359;
   wire n_5_1871;
   wire n_5_996;
   wire n_5_997;
   wire n_5_3360;
   wire n_5_998;
   wire n_5_999;
   wire n_5_2699;
   wire n_5_1000;
   wire n_5_1001;
   wire n_5_1002;
   wire n_5_1003;
   wire n_5_1004;
   wire n_5_1005;
   wire n_5_1923;
   wire n_5_1007;
   wire n_5_1008;
   wire n_5_1009;
   wire n_5_1010;
   wire n_5_1011;
   wire n_5_3364;
   wire n_5_1012;
   wire n_5_1013;
   wire n_5_3365;
   wire n_5_3366;
   wire n_5_3367;
   wire n_5_1014;
   wire n_5_1015;
   wire n_5_1924;
   wire n_5_1016;
   wire n_5_1017;
   wire n_5_1018;
   wire n_5_1019;
   wire n_5_1020;
   wire n_5_1021;
   wire n_5_1022;
   wire n_5_1023;
   wire n_5_3372;
   wire n_5_1024;
   wire n_5_1025;
   wire n_5_1026;
   wire n_5_1027;
   wire n_5_1028;
   wire n_5_1029;
   wire n_5_1030;
   wire n_5_456;
   wire n_5_460;
   wire n_5_4059;
   wire n_5_4060;
   wire n_5_4061;
   wire n_5_1033;
   wire n_5_1034;
   wire n_5_3377;
   wire n_5_1035;
   wire n_5_1036;
   wire n_5_1037;
   wire n_5_1038;
   wire n_5_1039;
   wire n_5_1938;
   wire n_5_1040;
   wire n_5_1041;
   wire n_5_1042;
   wire n_5_1043;
   wire n_5_1044;
   wire n_5_1045;
   wire n_5_1046;
   wire n_5_1047;
   wire n_5_1048;
   wire n_5_1049;
   wire n_5_1050;
   wire n_5_1051;
   wire n_5_4062;
   wire n_5_4063;
   wire n_5_1052;
   wire n_5_1053;
   wire n_5_1054;
   wire n_5_1055;
   wire n_5_1056;
   wire n_5_1057;
   wire n_5_1058;
   wire n_5_1059;
   wire n_5_1060;
   wire n_5_1061;
   wire n_5_1062;
   wire n_5_1063;
   wire n_5_1064;
   wire n_5_1065;
   wire n_5_1066;
   wire n_5_1067;
   wire n_5_1068;
   wire n_5_1069;
   wire n_5_1070;
   wire n_5_1071;
   wire n_5_1072;
   wire n_5_1073;
   wire n_5_3157;
   wire n_5_1074;
   wire n_5_1942;
   wire n_5_1075;
   wire n_5_4064;
   wire n_5_1076;
   wire n_5_1943;
   wire n_5_1077;
   wire n_5_1078;
   wire n_5_1079;
   wire n_5_1080;
   wire n_5_1081;
   wire n_5_1082;
   wire n_5_1083;
   wire n_5_1084;
   wire n_5_1085;
   wire n_5_1086;
   wire n_5_1087;
   wire n_5_1088;
   wire n_5_1089;
   wire n_5_1090;
   wire n_5_1091;
   wire n_5_1092;
   wire n_5_1093;
   wire n_5_1094;
   wire n_5_1095;
   wire n_5_1096;
   wire n_5_1097;
   wire n_5_1098;
   wire n_5_1099;
   wire n_5_1100;
   wire n_5_3158;
   wire n_5_1101;
   wire n_5_1102;
   wire n_5_1944;
   wire n_5_1103;
   wire n_5_1104;
   wire n_5_1105;
   wire n_5_1106;
   wire n_5_1107;
   wire n_5_1108;
   wire n_5_1109;
   wire n_5_1945;
   wire n_5_1110;
   wire n_5_1953;
   wire n_5_3379;
   wire n_5_3380;
   wire n_5_1111;
   wire n_5_1112;
   wire n_5_1113;
   wire n_5_1114;
   wire n_5_1115;
   wire n_5_1116;
   wire n_5_1117;
   wire n_5_1118;
   wire n_5_1119;
   wire n_5_1120;
   wire n_5_1121;
   wire n_5_1956;
   wire n_5_1122;
   wire n_5_1960;
   wire n_5_3381;
   wire n_5_1123;
   wire n_5_1124;
   wire n_5_1125;
   wire n_5_1126;
   wire n_5_1127;
   wire n_5_3160;
   wire n_5_3864;
   wire n_5_1128;
   wire n_5_3383;
   wire n_5_1962;
   wire n_5_1129;
   wire n_5_1968;
   wire n_5_1976;
   wire n_5_1978;
   wire n_5_1981;
   wire n_5_1130;
   wire n_5_1996;
   wire n_5_1131;
   wire n_5_1997;
   wire n_5_1132;
   wire n_5_1998;
   wire n_5_1133;
   wire n_5_1134;
   wire n_5_1135;
   wire n_5_1136;
   wire n_5_1137;
   wire n_5_1138;
   wire n_5_1139;
   wire n_5_1140;
   wire n_5_1141;
   wire n_5_1142;
   wire n_5_1143;
   wire n_5_1144;
   wire n_5_1145;
   wire n_5_1146;
   wire n_5_1147;
   wire n_5_1148;
   wire n_5_1149;
   wire n_5_1150;
   wire n_5_1151;
   wire n_5_1152;
   wire n_5_1153;
   wire n_5_1154;
   wire n_5_1999;
   wire n_5_2005;
   wire n_5_1155;
   wire n_5_1156;
   wire n_5_1157;
   wire n_5_1158;
   wire n_5_1159;
   wire n_5_1160;
   wire n_5_1161;
   wire n_5_1162;
   wire n_5_1163;
   wire n_5_1164;
   wire n_5_1165;
   wire n_5_1166;
   wire n_5_1167;
   wire n_5_1168;
   wire n_5_1169;
   wire n_5_2008;
   wire n_5_1170;
   wire n_5_1171;
   wire n_5_1172;
   wire n_5_1173;
   wire n_5_1174;
   wire n_5_1175;
   wire n_5_1176;
   wire n_5_1177;
   wire n_5_1178;
   wire n_5_1179;
   wire n_5_1180;
   wire n_5_1181;
   wire n_5_1182;
   wire n_5_1183;
   wire n_5_1184;
   wire n_5_1185;
   wire n_5_2016;
   wire n_5_1186;
   wire n_5_1187;
   wire n_5_1188;
   wire n_5_1189;
   wire n_5_1190;
   wire n_5_1191;
   wire n_5_1192;
   wire n_5_1193;
   wire n_5_1194;
   wire n_5_2023;
   wire n_5_1195;
   wire n_5_1196;
   wire n_5_2024;
   wire n_5_1197;
   wire n_5_2028;
   wire n_5_2029;
   wire n_5_1198;
   wire n_5_1199;
   wire n_5_2031;
   wire n_5_2032;
   wire n_5_1200;
   wire n_5_1201;
   wire n_5_1202;
   wire n_5_1203;
   wire n_5_1204;
   wire n_5_1205;
   wire n_5_1206;
   wire n_5_1207;
   wire n_5_1208;
   wire n_5_1209;
   wire n_5_1210;
   wire n_5_1211;
   wire n_5_2049;
   wire n_5_2050;
   wire n_5_2051;
   wire n_5_2088;
   wire n_5_2089;
   wire n_5_2090;
   wire n_5_2110;
   wire n_5_1212;
   wire n_5_3384;
   wire n_5_1213;
   wire n_5_2116;
   wire n_5_2153;
   wire n_5_2154;
   wire n_5_2155;
   wire n_5_2156;
   wire n_5_2157;
   wire n_5_2158;
   wire n_5_2159;
   wire n_5_2160;
   wire n_5_2161;
   wire n_5_2162;
   wire n_5_1214;
   wire n_5_3385;
   wire n_5_1215;
   wire n_5_1216;
   wire n_5_3386;
   wire n_5_1217;
   wire n_5_2165;
   wire n_5_2166;
   wire n_5_2167;
   wire n_5_1218;
   wire n_5_1219;
   wire n_5_1220;
   wire n_5_1221;
   wire n_5_1222;
   wire n_5_1223;
   wire n_5_1224;
   wire n_5_1946;
   wire n_5_1225;
   wire n_5_1226;
   wire n_5_1227;
   wire n_5_1228;
   wire n_5_1229;
   wire n_5_1230;
   wire n_5_1231;
   wire n_5_1232;
   wire n_5_1947;
   wire n_5_1950;
   wire n_5_1233;
   wire n_5_1234;
   wire n_5_1235;
   wire n_5_1236;
   wire n_5_1951;
   wire n_5_1237;
   wire n_5_1238;
   wire n_5_1239;
   wire n_5_1952;
   wire n_5_1240;
   wire n_5_1241;
   wire n_5_1242;
   wire n_5_1243;
   wire n_5_1954;
   wire n_5_1244;
   wire n_5_1245;
   wire n_5_1246;
   wire n_5_2168;
   wire n_5_1247;
   wire n_5_1248;
   wire n_5_2169;
   wire n_5_1249;
   wire n_5_1250;
   wire n_5_1251;
   wire n_5_1252;
   wire n_5_1253;
   wire n_5_1254;
   wire n_5_1255;
   wire n_5_1256;
   wire n_5_1257;
   wire n_5_2170;
   wire n_5_1258;
   wire n_5_1259;
   wire n_5_1260;
   wire n_5_1261;
   wire n_5_1262;
   wire n_5_1263;
   wire n_5_1264;
   wire n_5_1265;
   wire n_5_1266;
   wire n_5_1267;
   wire n_5_1268;
   wire n_5_1269;
   wire n_5_1270;
   wire n_5_1271;
   wire n_5_1272;
   wire n_5_1273;
   wire n_5_1274;
   wire n_5_1275;
   wire n_5_1276;
   wire n_5_1277;
   wire n_5_1278;
   wire n_5_1279;
   wire n_5_1280;
   wire n_5_1281;
   wire n_5_1282;
   wire n_5_1283;
   wire n_5_1284;
   wire n_5_1285;
   wire n_5_1286;
   wire n_5_1287;
   wire n_5_1288;
   wire n_5_1289;
   wire n_5_1290;
   wire n_5_1291;
   wire n_5_1292;
   wire n_5_1958;
   wire n_5_1293;
   wire n_5_1294;
   wire n_5_1295;
   wire n_5_1296;
   wire n_5_1297;
   wire n_5_1298;
   wire n_5_1959;
   wire n_5_1299;
   wire n_5_1803;
   wire n_5_1300;
   wire n_5_1301;
   wire n_5_1302;
   wire n_5_3162;
   wire n_5_1303;
   wire n_5_1304;
   wire n_5_1305;
   wire n_5_1306;
   wire n_5_1307;
   wire n_5_2174;
   wire n_5_1308;
   wire n_5_1309;
   wire n_5_1310;
   wire n_5_1311;
   wire n_5_1312;
   wire n_5_1313;
   wire n_5_1314;
   wire n_5_1315;
   wire n_5_1316;
   wire n_5_1317;
   wire n_5_1318;
   wire n_5_1319;
   wire n_5_1320;
   wire n_5_1321;
   wire n_5_1322;
   wire n_5_1323;
   wire n_5_1324;
   wire n_5_3163;
   wire n_5_1325;
   wire n_5_1326;
   wire n_5_2178;
   wire n_5_1327;
   wire n_5_1328;
   wire n_5_1329;
   wire n_5_1330;
   wire n_5_3164;
   wire n_5_1331;
   wire n_5_1332;
   wire n_5_1333;
   wire n_5_1334;
   wire n_5_1335;
   wire n_5_1336;
   wire n_5_1964;
   wire n_5_1337;
   wire n_5_1338;
   wire n_5_1339;
   wire n_5_1340;
   wire n_5_1341;
   wire n_5_1342;
   wire n_5_1966;
   wire n_5_1967;
   wire n_5_2179;
   wire n_5_2180;
   wire n_5_2181;
   wire n_5_1343;
   wire n_5_1969;
   wire n_5_1970;
   wire n_5_3165;
   wire n_5_3166;
   wire n_5_3167;
   wire n_5_1344;
   wire n_5_1345;
   wire n_5_1971;
   wire n_5_1346;
   wire n_5_1347;
   wire n_5_1348;
   wire n_5_1349;
   wire n_5_1350;
   wire n_5_1351;
   wire n_5_1352;
   wire n_5_1353;
   wire n_5_1354;
   wire n_5_1355;
   wire n_5_1356;
   wire n_5_1357;
   wire n_5_1358;
   wire n_5_2182;
   wire n_5_1359;
   wire n_5_1360;
   wire n_5_1361;
   wire n_5_1362;
   wire n_5_1363;
   wire n_5_1364;
   wire n_5_1365;
   wire n_5_1366;
   wire n_5_1367;
   wire n_5_1368;
   wire n_5_1369;
   wire n_5_1370;
   wire n_5_1371;
   wire n_5_1372;
   wire n_5_461;
   wire n_5_1375;
   wire n_5_1376;
   wire n_5_1377;
   wire n_5_1378;
   wire n_5_1972;
   wire n_5_1379;
   wire n_5_1973;
   wire n_5_1380;
   wire n_5_1974;
   wire n_5_3387;
   wire n_5_1381;
   wire n_5_1977;
   wire n_5_1979;
   wire n_5_1383;
   wire n_5_1384;
   wire n_5_1385;
   wire n_5_2185;
   wire n_5_1386;
   wire n_5_1387;
   wire n_5_1980;
   wire n_5_1388;
   wire n_5_1389;
   wire n_5_1390;
   wire n_5_2186;
   wire n_5_1982;
   wire n_5_1983;
   wire n_5_1391;
   wire n_5_1392;
   wire n_5_2187;
   wire n_5_1393;
   wire n_5_2188;
   wire n_5_1394;
   wire n_5_1395;
   wire n_5_1984;
   wire n_5_1396;
   wire n_5_1397;
   wire n_5_1398;
   wire n_5_1399;
   wire n_5_1400;
   wire n_5_1401;
   wire n_5_1402;
   wire n_5_1403;
   wire n_5_1404;
   wire n_5_1405;
   wire n_5_1406;
   wire n_5_1407;
   wire n_5_1408;
   wire n_5_2189;
   wire n_5_1409;
   wire n_5_1410;
   wire n_5_1411;
   wire n_5_1412;
   wire n_5_1413;
   wire n_5_2190;
   wire n_5_1414;
   wire n_5_1986;
   wire n_5_1415;
   wire n_5_1987;
   wire n_5_1416;
   wire n_5_1417;
   wire n_5_1418;
   wire n_5_1419;
   wire n_5_1420;
   wire n_5_1421;
   wire n_5_1988;
   wire n_5_1422;
   wire n_5_1423;
   wire n_5_1989;
   wire n_5_1424;
   wire n_5_1425;
   wire n_5_1426;
   wire n_5_1427;
   wire n_5_1428;
   wire n_5_1429;
   wire n_5_1430;
   wire n_5_1431;
   wire n_5_1432;
   wire n_5_1433;
   wire n_5_1434;
   wire n_5_1435;
   wire n_5_1436;
   wire n_5_1437;
   wire n_5_1438;
   wire n_5_1439;
   wire n_5_2191;
   wire n_5_2192;
   wire n_5_1440;
   wire n_5_1441;
   wire n_5_3168;
   wire n_5_1442;
   wire n_5_1443;
   wire n_5_1444;
   wire n_5_1445;
   wire n_5_1446;
   wire n_5_1447;
   wire n_5_1448;
   wire n_5_1449;
   wire n_5_1450;
   wire n_5_1451;
   wire n_5_1452;
   wire n_5_3170;
   wire n_5_1453;
   wire n_5_3171;
   wire n_5_1454;
   wire n_5_2196;
   wire n_5_1455;
   wire n_5_1456;
   wire n_5_1457;
   wire n_5_2197;
   wire n_5_2198;
   wire n_5_2199;
   wire n_5_3172;
   wire n_5_4065;
   wire n_5_1458;
   wire n_5_1459;
   wire n_5_1460;
   wire n_5_1461;
   wire n_5_3173;
   wire n_5_3174;
   wire n_5_2202;
   wire n_5_1462;
   wire n_5_1463;
   wire n_5_1464;
   wire n_5_1465;
   wire n_5_1466;
   wire n_5_1467;
   wire n_5_1468;
   wire n_5_2203;
   wire n_5_1469;
   wire n_5_1470;
   wire n_5_2204;
   wire n_5_2206;
   wire n_5_1471;
   wire n_5_3175;
   wire n_5_1472;
   wire n_5_1473;
   wire n_5_3176;
   wire n_5_1474;
   wire n_5_1475;
   wire n_5_1476;
   wire n_5_2000;
   wire n_5_1477;
   wire n_5_1478;
   wire n_5_1479;
   wire n_5_2001;
   wire n_5_1480;
   wire n_5_2207;
   wire n_5_1481;
   wire n_5_1482;
   wire n_5_1483;
   wire n_5_2208;
   wire n_5_1484;
   wire n_5_2209;
   wire n_5_1485;
   wire n_5_1486;
   wire n_5_1487;
   wire n_5_1488;
   wire n_5_1489;
   wire n_5_1490;
   wire n_5_1491;
   wire n_5_1492;
   wire n_5_1493;
   wire n_5_1494;
   wire n_5_1495;
   wire n_5_1496;
   wire n_5_1497;
   wire n_5_1498;
   wire n_5_1499;
   wire n_5_2210;
   wire n_5_1500;
   wire n_5_1501;
   wire n_5_1502;
   wire n_5_1804;
   wire n_5_1503;
   wire n_5_1504;
   wire n_5_1505;
   wire n_5_1506;
   wire n_5_1507;
   wire n_5_1508;
   wire n_5_1509;
   wire n_5_3177;
   wire n_5_1510;
   wire n_5_1511;
   wire n_5_1512;
   wire n_5_1513;
   wire n_5_1514;
   wire n_5_1515;
   wire n_5_1516;
   wire n_5_1517;
   wire n_5_1518;
   wire n_5_1519;
   wire n_5_1520;
   wire n_5_1521;
   wire n_5_2002;
   wire n_5_2003;
   wire n_5_1522;
   wire n_5_1523;
   wire n_5_1524;
   wire n_5_1525;
   wire n_5_1526;
   wire n_5_1527;
   wire n_5_1528;
   wire n_5_1529;
   wire n_5_1530;
   wire n_5_1531;
   wire n_5_1532;
   wire n_5_1533;
   wire n_5_1534;
   wire n_5_1535;
   wire n_5_1536;
   wire n_5_1537;
   wire n_5_1538;
   wire n_5_1539;
   wire n_5_1540;
   wire n_5_1541;
   wire n_5_1542;
   wire n_5_1543;
   wire n_5_1544;
   wire n_5_1545;
   wire n_5_1546;
   wire n_5_1547;
   wire n_5_1548;
   wire n_5_1549;
   wire n_5_2004;
   wire n_5_1550;
   wire n_5_1551;
   wire n_5_2211;
   wire n_5_1552;
   wire n_5_1553;
   wire n_5_2212;
   wire n_5_1554;
   wire n_5_2213;
   wire n_5_1555;
   wire n_5_1556;
   wire n_5_1557;
   wire n_5_1558;
   wire n_5_1559;
   wire n_5_1560;
   wire n_5_1561;
   wire n_5_1562;
   wire n_5_1563;
   wire n_5_2006;
   wire n_5_1564;
   wire n_5_1565;
   wire n_5_1566;
   wire n_5_1567;
   wire n_5_1568;
   wire n_5_1569;
   wire n_5_1570;
   wire n_5_1571;
   wire n_5_1572;
   wire n_5_2007;
   wire n_5_1573;
   wire n_5_1574;
   wire n_5_1575;
   wire n_5_1576;
   wire n_5_1577;
   wire n_5_1578;
   wire n_5_1579;
   wire n_5_1580;
   wire n_5_1581;
   wire n_5_1582;
   wire n_5_1583;
   wire n_5_1805;
   wire n_5_1584;
   wire n_5_1585;
   wire n_5_1586;
   wire n_5_1587;
   wire n_5_1588;
   wire n_5_1589;
   wire n_5_2214;
   wire n_5_1590;
   wire n_5_1591;
   wire n_5_1592;
   wire n_5_1593;
   wire n_5_1594;
   wire n_5_3178;
   wire n_5_2216;
   wire n_5_1595;
   wire n_5_1596;
   wire n_5_1597;
   wire n_5_1598;
   wire n_5_1599;
   wire n_5_1600;
   wire n_5_1601;
   wire n_5_1602;
   wire n_5_1603;
   wire n_5_1604;
   wire n_5_1605;
   wire n_5_1606;
   wire n_5_2217;
   wire n_5_1607;
   wire n_5_1608;
   wire n_5_1609;
   wire n_5_1610;
   wire n_5_1611;
   wire n_5_1612;
   wire n_5_1613;
   wire n_5_1614;
   wire n_5_1615;
   wire n_5_1616;
   wire n_5_1617;
   wire n_5_1618;
   wire n_5_1619;
   wire n_5_1620;
   wire n_5_1621;
   wire n_5_2218;
   wire n_5_1622;
   wire n_5_2219;
   wire n_5_1623;
   wire n_5_1624;
   wire n_5_1625;
   wire n_5_1626;
   wire n_5_1627;
   wire n_5_1628;
   wire n_5_1629;
   wire n_5_1630;
   wire n_5_1631;
   wire n_5_1632;
   wire n_5_1633;
   wire n_5_1634;
   wire n_5_1635;
   wire n_5_1636;
   wire n_5_1637;
   wire n_5_1638;
   wire n_5_1639;
   wire n_5_1640;
   wire n_5_1641;
   wire n_5_1642;
   wire n_5_1643;
   wire n_5_1644;
   wire n_5_1645;
   wire n_5_1646;
   wire n_5_1647;
   wire n_5_1648;
   wire n_5_1649;
   wire n_5_1650;
   wire n_5_1651;
   wire n_5_1652;
   wire n_5_1653;
   wire n_5_1654;
   wire n_5_1655;
   wire n_5_1656;
   wire n_5_1657;
   wire n_5_3179;
   wire n_5_1658;
   wire n_5_1659;
   wire n_5_1660;
   wire n_5_1661;
   wire n_5_1662;
   wire n_5_1663;
   wire n_5_1664;
   wire n_5_1665;
   wire n_5_1666;
   wire n_5_1667;
   wire n_5_1668;
   wire n_5_1669;
   wire n_5_1670;
   wire n_5_1671;
   wire n_5_1672;
   wire n_5_1673;
   wire n_5_1674;
   wire n_5_1675;
   wire n_5_1676;
   wire n_5_1677;
   wire n_5_1678;
   wire n_5_1679;
   wire n_5_1680;
   wire n_5_1681;
   wire n_5_1682;
   wire n_5_1683;
   wire n_5_1684;
   wire n_5_1685;
   wire n_5_4066;
   wire n_5_1686;
   wire n_5_1687;
   wire n_5_1688;
   wire n_5_1689;
   wire n_5_1690;
   wire n_5_1691;
   wire n_5_1692;
   wire n_5_1693;
   wire n_5_1694;
   wire n_5_1695;
   wire n_5_1696;
   wire n_5_1697;
   wire n_5_1698;
   wire n_5_1699;
   wire n_5_2221;
   wire n_5_1700;
   wire n_5_1701;
   wire n_5_1702;
   wire n_5_1703;
   wire n_5_1704;
   wire n_5_1705;
   wire n_5_1706;
   wire n_5_1707;
   wire n_5_1708;
   wire n_5_1709;
   wire n_5_1710;
   wire n_5_1711;
   wire n_5_3180;
   wire n_5_3181;
   wire n_5_1712;
   wire n_5_1713;
   wire n_5_1714;
   wire n_5_1715;
   wire n_5_1716;
   wire n_5_1717;
   wire n_5_1718;
   wire n_5_1719;
   wire n_5_1720;
   wire n_5_1721;
   wire n_5_2225;
   wire n_5_1722;
   wire n_5_1723;
   wire n_5_2010;
   wire n_5_2011;
   wire n_5_1724;
   wire n_5_2012;
   wire n_5_1725;
   wire n_5_1726;
   wire n_5_1727;
   wire n_5_1728;
   wire n_5_1729;
   wire n_5_1730;
   wire n_5_1731;
   wire n_5_1732;
   wire n_5_1733;
   wire n_5_3182;
   wire n_5_1734;
   wire n_5_2013;
   wire n_5_1735;
   wire n_5_1736;
   wire n_5_1737;
   wire n_5_1738;
   wire n_5_1739;
   wire n_5_1740;
   wire n_5_1741;
   wire n_5_1742;
   wire n_5_1743;
   wire n_5_1744;
   wire n_5_1745;
   wire n_5_1746;
   wire n_5_1747;
   wire n_5_1748;
   wire n_5_2014;
   wire n_5_1749;
   wire n_5_1750;
   wire n_5_1751;
   wire n_5_1752;
   wire n_5_1753;
   wire n_5_1754;
   wire n_5_2228;
   wire n_5_1755;
   wire n_5_1756;
   wire n_5_1808;
   wire n_5_1810;
   wire n_5_1757;
   wire n_5_1758;
   wire n_5_1759;
   wire n_5_1760;
   wire n_5_1761;
   wire n_5_1762;
   wire n_5_3183;
   wire n_5_1763;
   wire n_5_1764;
   wire n_5_1765;
   wire n_5_1766;
   wire n_5_1767;
   wire n_5_1768;
   wire n_5_1769;
   wire n_5_1770;
   wire n_5_2017;
   wire n_5_2229;
   wire n_5_1771;
   wire n_5_1772;
   wire n_5_1773;
   wire n_5_1774;
   wire n_5_1775;
   wire n_5_1776;
   wire n_5_1777;
   wire n_5_1778;
   wire n_5_1779;
   wire n_5_1780;
   wire n_5_1781;
   wire n_5_1782;
   wire n_5_1783;
   wire n_5_1784;
   wire n_5_1785;
   wire n_5_1786;
   wire n_5_1787;
   wire n_5_1790;
   wire n_5_1788;
   wire n_5_1789;
   wire n_5_1791;
   wire n_5_1792;
   wire n_5_2022;
   wire n_5_2232;
   wire n_5_2233;
   wire n_5_2234;
   wire n_5_2025;
   wire n_5_2235;
   wire n_5_2236;
   wire n_5_2237;
   wire n_5_1793;
   wire n_5_1794;
   wire n_5_1795;
   wire n_5_1811;
   wire n_5_1796;
   wire n_5_1797;
   wire n_5_1798;
   wire n_5_1812;
   wire n_5_1799;
   wire n_5_1813;
   wire n_5_2238;
   wire n_5_1800;
   wire n_5_2239;
   wire n_5_1801;
   wire n_5_3389;
   wire n_5_1802;
   wire n_5_1807;
   wire n_5_1809;
   wire n_5_1816;
   wire n_5_2240;
   wire n_5_2241;
   wire n_5_2242;
   wire n_5_2243;
   wire n_5_4067;
   wire n_5_1814;
   wire n_5_1815;
   wire n_5_1818;
   wire n_5_1821;
   wire n_5_1822;
   wire n_5_1823;
   wire n_5_4068;
   wire n_5_2245;
   wire n_5_4069;
   wire n_5_2247;
   wire n_5_1824;
   wire n_5_2248;
   wire n_5_1825;
   wire n_5_1827;
   wire n_5_1829;
   wire n_5_1830;
   wire n_5_2249;
   wire n_5_2250;
   wire n_5_2251;
   wire n_5_2252;
   wire n_5_1831;
   wire n_5_1832;
   wire n_5_1833;
   wire n_5_1834;
   wire n_5_1835;
   wire n_5_1836;
   wire n_5_1837;
   wire n_5_1838;
   wire n_5_1839;
   wire n_5_1840;
   wire n_5_1841;
   wire n_5_1842;
   wire n_5_1843;
   wire n_5_1845;
   wire n_5_1846;
   wire n_5_1847;
   wire n_5_1848;
   wire n_5_1849;
   wire n_5_1851;
   wire n_5_1852;
   wire n_5_1853;
   wire n_5_1854;
   wire n_5_2253;
   wire n_5_1855;
   wire n_5_1856;
   wire n_5_1857;
   wire n_5_1858;
   wire n_5_1859;
   wire n_5_1860;
   wire n_5_1861;
   wire n_5_1862;
   wire n_5_1864;
   wire n_5_1865;
   wire n_5_1866;
   wire n_5_3392;
   wire n_5_1867;
   wire n_5_1868;
   wire n_5_1869;
   wire n_5_1870;
   wire n_5_1872;
   wire n_5_1873;
   wire n_5_1874;
   wire n_5_1875;
   wire n_5_1876;
   wire n_5_1877;
   wire n_5_1878;
   wire n_5_1879;
   wire n_5_1880;
   wire n_5_1881;
   wire n_5_1882;
   wire n_5_1883;
   wire n_5_1884;
   wire n_5_1885;
   wire n_5_1886;
   wire n_5_1887;
   wire n_5_1888;
   wire n_5_1889;
   wire n_5_2254;
   wire n_5_1890;
   wire n_5_2255;
   wire n_5_1891;
   wire n_5_1892;
   wire n_5_1893;
   wire n_5_4070;
   wire n_5_1894;
   wire n_5_1895;
   wire n_5_1896;
   wire n_5_1897;
   wire n_5_2256;
   wire n_5_1898;
   wire n_5_1899;
   wire n_5_1900;
   wire n_5_1901;
   wire n_5_1902;
   wire n_5_1903;
   wire n_5_1904;
   wire n_5_1905;
   wire n_5_1906;
   wire n_5_1907;
   wire n_5_1908;
   wire n_5_1909;
   wire n_5_1910;
   wire n_5_1911;
   wire n_5_1912;
   wire n_5_1913;
   wire n_5_1914;
   wire n_5_1915;
   wire n_5_1916;
   wire n_5_1917;
   wire n_5_1918;
   wire n_5_1919;
   wire n_5_1920;
   wire n_5_1921;
   wire n_5_1922;
   wire n_5_1925;
   wire n_5_1926;
   wire n_5_1927;
   wire n_5_1928;
   wire n_5_1929;
   wire n_5_1930;
   wire n_5_1931;
   wire n_5_1932;
   wire n_5_1933;
   wire n_5_1934;
   wire n_5_1935;
   wire n_5_1936;
   wire n_5_1937;
   wire n_5_1939;
   wire n_5_1940;
   wire n_5_1941;
   wire n_5_1948;
   wire n_5_1949;
   wire n_5_1955;
   wire n_5_1957;
   wire n_5_1961;
   wire n_5_1963;
   wire n_5_1965;
   wire n_5_2257;
   wire n_5_2258;
   wire n_5_1975;
   wire n_5_1985;
   wire n_5_1990;
   wire n_5_1991;
   wire n_5_1992;
   wire n_5_1993;
   wire n_5_1994;
   wire n_5_2259;
   wire n_5_1995;
   wire n_5_2260;
   wire n_5_2009;
   wire n_5_2015;
   wire n_5_2018;
   wire n_5_2019;
   wire n_5_2020;
   wire n_5_2021;
   wire n_5_2026;
   wire n_5_2027;
   wire n_5_2030;
   wire n_5_2033;
   wire n_5_2034;
   wire n_5_2035;
   wire n_5_2036;
   wire n_5_2037;
   wire n_5_2038;
   wire n_5_2039;
   wire n_5_2040;
   wire n_5_2041;
   wire n_5_2042;
   wire n_5_2043;
   wire n_5_2044;
   wire n_5_2045;
   wire n_5_2046;
   wire n_5_2047;
   wire n_5_2048;
   wire n_5_2052;
   wire n_5_2053;
   wire n_5_2054;
   wire n_5_2055;
   wire n_5_2056;
   wire n_5_2057;
   wire n_5_2058;
   wire n_5_2059;
   wire n_5_2060;
   wire n_5_2061;
   wire n_5_2062;
   wire n_5_2063;
   wire n_5_2064;
   wire n_5_2065;
   wire n_5_2066;
   wire n_5_2067;
   wire n_5_2068;
   wire n_5_2069;
   wire n_5_2070;
   wire n_5_2071;
   wire n_5_2072;
   wire n_5_2073;
   wire n_5_2261;
   wire n_5_2074;
   wire n_5_2075;
   wire n_5_2076;
   wire n_5_2077;
   wire n_5_2078;
   wire n_5_2079;
   wire n_5_2080;
   wire n_5_2081;
   wire n_5_2082;
   wire n_5_2083;
   wire n_5_2084;
   wire n_5_2085;
   wire n_5_2086;
   wire n_5_2087;
   wire n_5_2091;
   wire n_5_2092;
   wire n_5_2093;
   wire n_5_2094;
   wire n_5_2095;
   wire n_5_2096;
   wire n_5_2097;
   wire n_5_2098;
   wire n_5_2099;
   wire n_5_2100;
   wire n_5_2101;
   wire n_5_2102;
   wire n_5_2103;
   wire n_5_2104;
   wire n_5_2105;
   wire n_5_2106;
   wire n_5_2107;
   wire n_5_2108;
   wire n_5_2109;
   wire n_5_2111;
   wire n_5_2112;
   wire n_5_2113;
   wire n_5_2114;
   wire n_5_2115;
   wire n_5_2117;
   wire n_5_2262;
   wire n_5_2118;
   wire n_5_2119;
   wire n_5_2120;
   wire n_5_2121;
   wire n_5_2122;
   wire n_5_2123;
   wire n_5_2263;
   wire n_5_2124;
   wire n_5_2264;
   wire n_5_2265;
   wire n_5_2125;
   wire n_5_2266;
   wire n_5_2126;
   wire n_5_3393;
   wire n_5_2127;
   wire n_5_2267;
   wire n_5_2128;
   wire n_5_2129;
   wire n_5_4071;
   wire n_5_2130;
   wire n_5_2268;
   wire n_5_2131;
   wire n_5_2132;
   wire n_5_2133;
   wire n_5_2134;
   wire n_5_2135;
   wire n_5_2136;
   wire n_5_2137;
   wire n_5_2138;
   wire n_5_2139;
   wire n_5_2269;
   wire n_5_2140;
   wire n_5_2141;
   wire n_5_2142;
   wire n_5_2143;
   wire n_5_2144;
   wire n_5_2145;
   wire n_5_2146;
   wire n_5_2147;
   wire n_5_2148;
   wire n_5_2149;
   wire n_5_2150;
   wire n_5_2151;
   wire n_5_2152;
   wire n_5_2163;
   wire n_5_2164;
   wire n_5_2171;
   wire n_5_2172;
   wire n_5_2173;
   wire n_5_2175;
   wire n_5_2176;
   wire n_5_2177;
   wire n_5_2183;
   wire n_5_2193;
   wire n_5_2194;
   wire n_5_2195;
   wire n_5_2200;
   wire n_5_2201;
   wire n_5_2270;
   wire n_5_2205;
   wire n_5_2215;
   wire n_5_2220;
   wire n_5_2222;
   wire n_5_2223;
   wire n_5_2224;
   wire n_5_2226;
   wire n_5_2227;
   wire n_5_2230;
   wire n_5_2231;
   wire n_5_2244;
   wire n_5_2271;
   wire n_5_2246;
   wire n_5_2272;
   wire n_5_2273;
   wire n_5_2274;
   wire n_5_2275;
   wire n_5_2276;
   wire n_5_2277;
   wire n_5_2278;
   wire n_5_2279;
   wire n_5_2280;
   wire n_5_2281;
   wire n_5_2282;
   wire n_5_2283;
   wire n_5_2284;
   wire n_5_2285;
   wire n_5_2286;
   wire n_5_2287;
   wire n_5_2288;
   wire n_5_2289;
   wire n_5_2290;
   wire n_5_2291;
   wire n_5_2292;
   wire n_5_2293;
   wire n_5_2294;
   wire n_5_2295;
   wire n_5_2296;
   wire n_5_2297;
   wire n_5_2298;
   wire n_5_2299;
   wire n_5_2300;
   wire n_5_2301;
   wire n_5_2302;
   wire n_5_2303;
   wire n_5_2304;
   wire n_5_2305;
   wire n_5_2306;
   wire n_5_2307;
   wire n_5_2308;
   wire n_5_2309;
   wire n_5_2310;
   wire n_5_2311;
   wire n_5_2312;
   wire n_5_2313;
   wire n_5_2314;
   wire n_5_2315;
   wire n_5_2316;
   wire n_5_2317;
   wire n_5_2318;
   wire n_5_2319;
   wire n_5_2320;
   wire n_5_2321;
   wire n_5_2322;
   wire n_5_2323;
   wire n_5_2324;
   wire n_5_2325;
   wire n_5_2326;
   wire n_5_2327;
   wire n_5_2328;
   wire n_5_2329;
   wire n_5_2330;
   wire n_5_2331;
   wire n_5_2332;
   wire n_5_2333;
   wire n_5_2334;
   wire n_5_2335;
   wire n_5_2336;
   wire n_5_2337;
   wire n_5_2338;
   wire n_5_2339;
   wire n_5_2340;
   wire n_5_2341;
   wire n_5_2342;
   wire n_5_2343;
   wire n_5_2344;
   wire n_5_2345;
   wire n_5_2346;
   wire n_5_2347;
   wire n_5_2348;
   wire n_5_4072;
   wire n_5_2349;
   wire n_5_2350;
   wire n_5_2351;
   wire n_5_2352;
   wire n_5_2353;
   wire n_5_2354;
   wire n_5_2355;
   wire n_5_2356;
   wire n_5_2357;
   wire n_5_2358;
   wire n_5_2359;
   wire n_5_2360;
   wire n_5_2361;
   wire n_5_2362;
   wire n_5_2363;
   wire n_5_2364;
   wire n_5_2365;
   wire n_5_2366;
   wire n_5_2367;
   wire n_5_2368;
   wire n_5_2369;
   wire n_5_2370;
   wire n_5_2371;
   wire n_5_2372;
   wire n_5_2373;
   wire n_5_2374;
   wire n_5_2375;
   wire n_5_2376;
   wire n_5_2377;
   wire n_5_2378;
   wire n_5_2379;
   wire n_5_2380;
   wire n_5_2381;
   wire n_5_2382;
   wire n_5_2383;
   wire n_5_2384;
   wire n_5_2385;
   wire n_5_2386;
   wire n_5_2387;
   wire n_5_2388;
   wire n_5_2389;
   wire n_5_2390;
   wire n_5_4073;
   wire n_5_2391;
   wire n_5_2392;
   wire n_5_2393;
   wire n_5_2394;
   wire n_5_2395;
   wire n_5_2396;
   wire n_5_2397;
   wire n_5_2398;
   wire n_5_2399;
   wire n_5_2400;
   wire n_5_2401;
   wire n_5_2402;
   wire n_5_2403;
   wire n_5_2404;
   wire n_5_2405;
   wire n_5_2406;
   wire n_5_2407;
   wire n_5_2408;
   wire n_5_2409;
   wire n_5_2410;
   wire n_5_2411;
   wire n_5_2412;
   wire n_5_2413;
   wire n_5_2414;
   wire n_5_2415;
   wire n_5_2416;
   wire n_5_2417;
   wire n_5_2418;
   wire n_5_2419;
   wire n_5_2420;
   wire n_5_2421;
   wire n_5_2422;
   wire n_5_2423;
   wire n_5_2424;
   wire n_5_2425;
   wire n_5_2426;
   wire n_5_2427;
   wire n_5_2428;
   wire n_5_2429;
   wire n_5_2430;
   wire n_5_2431;
   wire n_5_2432;
   wire n_5_2433;
   wire n_5_2434;
   wire n_5_2435;
   wire n_5_2436;
   wire n_5_2437;
   wire n_5_2438;
   wire n_5_2439;
   wire n_5_2440;
   wire n_5_2441;
   wire n_5_2442;
   wire n_5_2443;
   wire n_5_2444;
   wire n_5_2445;
   wire n_5_2446;
   wire n_5_2447;
   wire n_5_2448;
   wire n_5_2449;
   wire n_5_2450;
   wire n_5_2451;
   wire n_5_2452;
   wire n_5_2453;
   wire n_5_2454;
   wire n_5_2455;
   wire n_5_2456;
   wire n_5_2457;
   wire n_5_2458;
   wire n_5_2459;
   wire n_5_2460;
   wire n_5_2461;
   wire n_5_2462;
   wire n_5_2463;
   wire n_5_2464;
   wire n_5_2465;
   wire n_5_2466;
   wire n_5_2467;
   wire n_5_2468;
   wire n_5_2469;
   wire n_5_2470;
   wire n_5_2471;
   wire n_5_2472;
   wire n_5_2473;
   wire n_5_2474;
   wire n_5_2475;
   wire n_5_2476;
   wire n_5_2477;
   wire n_5_2478;
   wire n_5_2479;
   wire n_5_2480;
   wire n_5_2481;
   wire n_5_2482;
   wire n_5_2483;
   wire n_5_2484;
   wire n_5_2485;
   wire n_5_2486;
   wire n_5_2487;
   wire n_5_2488;
   wire n_5_2489;
   wire n_5_2490;
   wire n_5_2491;
   wire n_5_2492;
   wire n_5_2493;
   wire n_5_2494;
   wire n_5_2495;
   wire n_5_4074;
   wire n_5_2496;
   wire n_5_2497;
   wire n_5_2498;
   wire n_5_2499;
   wire n_5_2500;
   wire n_5_2501;
   wire n_5_2502;
   wire n_5_2503;
   wire n_5_2504;
   wire n_5_2505;
   wire n_5_2506;
   wire n_5_2507;
   wire n_5_2508;
   wire n_5_2509;
   wire n_5_2510;
   wire n_5_2511;
   wire n_5_2512;
   wire n_5_2513;
   wire n_5_4075;
   wire n_5_4076;
   wire n_5_4077;
   wire n_5_2514;
   wire n_5_2515;
   wire n_5_2516;
   wire n_5_2517;
   wire n_5_2518;
   wire n_5_2519;
   wire n_5_2520;
   wire n_5_2521;
   wire n_5_2522;
   wire n_5_2523;
   wire n_5_2524;
   wire n_5_2525;
   wire n_5_2526;
   wire n_5_2527;
   wire n_5_2528;
   wire n_5_2529;
   wire n_5_2530;
   wire n_5_2531;
   wire n_5_2532;
   wire n_5_2533;
   wire n_5_2534;
   wire n_5_2535;
   wire n_5_2536;
   wire n_5_2537;
   wire n_5_2538;
   wire n_5_2539;
   wire n_5_2540;
   wire n_5_2541;
   wire n_5_2542;
   wire n_5_2543;
   wire n_5_2544;
   wire n_5_2545;
   wire n_5_2546;
   wire n_5_2547;
   wire n_5_2548;
   wire n_5_2549;
   wire n_5_2550;
   wire n_5_2551;
   wire n_5_2552;
   wire n_5_2553;
   wire n_5_2554;
   wire n_5_2555;
   wire n_5_2556;
   wire n_5_2557;
   wire n_5_2558;
   wire n_5_2559;
   wire n_5_2560;
   wire n_5_2561;
   wire n_5_2562;
   wire n_5_2563;
   wire n_5_2564;
   wire n_5_2565;
   wire n_5_2566;
   wire n_5_2567;
   wire n_5_2568;
   wire n_5_2569;
   wire n_5_2570;
   wire n_5_2571;
   wire n_5_2572;
   wire n_5_2573;
   wire n_5_2574;
   wire n_5_2575;
   wire n_5_2576;
   wire n_5_2577;
   wire n_5_2578;
   wire n_5_2579;
   wire n_5_2580;
   wire n_5_2581;
   wire n_5_2582;
   wire n_5_2583;
   wire n_5_2584;
   wire n_5_2585;
   wire n_5_2586;
   wire n_5_2587;
   wire n_5_2588;
   wire n_5_2589;
   wire n_5_2590;
   wire n_5_2591;
   wire n_5_2592;
   wire n_5_2593;
   wire n_5_2594;
   wire n_5_2595;
   wire n_5_2596;
   wire n_5_2597;
   wire n_5_2598;
   wire n_5_3185;
   wire n_5_2599;
   wire n_5_2600;
   wire n_5_2601;
   wire n_5_2602;
   wire n_5_2603;
   wire n_5_2604;
   wire n_5_2605;
   wire n_5_2606;
   wire n_5_2607;
   wire n_5_2608;
   wire n_5_2609;
   wire n_5_2610;
   wire n_5_2611;
   wire n_5_2612;
   wire n_5_2613;
   wire n_5_2614;
   wire n_5_2615;
   wire n_5_2616;
   wire n_5_2617;
   wire n_5_2618;
   wire n_5_2619;
   wire n_5_2620;
   wire n_5_2621;
   wire n_5_2622;
   wire n_5_2623;
   wire n_5_2624;
   wire n_5_2625;
   wire n_5_2626;
   wire n_5_2627;
   wire n_5_2628;
   wire n_5_2629;
   wire n_5_2630;
   wire n_5_2631;
   wire n_5_2632;
   wire n_5_2633;
   wire n_5_2634;
   wire n_5_2635;
   wire n_5_2636;
   wire n_5_2637;
   wire n_5_2638;
   wire n_5_2639;
   wire n_5_2640;
   wire n_5_2641;
   wire n_5_2642;
   wire n_5_2643;
   wire n_5_2644;
   wire n_5_2645;
   wire n_5_2646;
   wire n_5_2647;
   wire n_5_2648;
   wire n_5_2649;
   wire n_5_2650;
   wire n_5_2651;
   wire n_5_2652;
   wire n_5_2653;
   wire n_5_2654;
   wire n_5_2655;
   wire n_5_2656;
   wire n_5_2657;
   wire n_5_2658;
   wire n_5_2659;
   wire n_5_2660;
   wire n_5_2661;
   wire n_5_2662;
   wire n_5_2663;
   wire n_5_2664;
   wire n_5_2665;
   wire n_5_2666;
   wire n_5_2667;
   wire n_5_2668;
   wire n_5_2669;
   wire n_5_2670;
   wire n_5_2671;
   wire n_5_2672;
   wire n_5_2673;
   wire n_5_2674;
   wire n_5_2675;
   wire n_5_2676;
   wire n_5_2677;
   wire n_5_2678;
   wire n_5_2679;
   wire n_5_2680;
   wire n_5_2681;
   wire n_5_2682;
   wire n_5_2683;
   wire n_5_2684;
   wire n_5_2685;
   wire n_5_2686;
   wire n_5_2687;
   wire n_5_2688;
   wire n_5_2689;
   wire n_5_2690;
   wire n_5_2691;
   wire n_5_2692;
   wire n_5_2693;
   wire n_5_2694;
   wire n_5_2695;
   wire n_5_2696;
   wire n_5_2697;
   wire n_5_2698;
   wire n_5_2700;
   wire n_5_2701;
   wire n_5_2702;
   wire n_5_2703;
   wire n_5_2704;
   wire n_5_2705;
   wire n_5_2706;
   wire n_5_2707;
   wire n_5_2708;
   wire n_5_2709;
   wire n_5_2710;
   wire n_5_2711;
   wire n_5_2712;
   wire n_5_2713;
   wire n_5_2714;
   wire n_5_2715;
   wire n_5_2716;
   wire n_5_2717;
   wire n_5_2718;
   wire n_5_2719;
   wire n_5_2720;
   wire n_5_2721;
   wire n_5_2722;
   wire n_5_2723;
   wire n_5_2724;
   wire n_5_2725;
   wire n_5_2726;
   wire n_5_2727;
   wire n_5_2728;
   wire n_5_2729;
   wire n_5_2730;
   wire n_5_2731;
   wire n_5_2732;
   wire n_5_2733;
   wire n_5_2734;
   wire n_5_2735;
   wire n_5_2736;
   wire n_5_2737;
   wire n_5_2738;
   wire n_5_2739;
   wire n_5_2740;
   wire n_5_2741;
   wire n_5_2742;
   wire n_5_2743;
   wire n_5_2744;
   wire n_5_2745;
   wire n_5_2746;
   wire n_5_2747;
   wire n_5_2748;
   wire n_5_2749;
   wire n_5_2750;
   wire n_5_2751;
   wire n_5_2752;
   wire n_5_2753;
   wire n_5_2754;
   wire n_5_2755;
   wire n_5_2756;
   wire n_5_2757;
   wire n_5_2758;
   wire n_5_2759;
   wire n_5_2760;
   wire n_5_2761;
   wire n_5_2762;
   wire n_5_2763;
   wire n_5_2764;
   wire n_5_2765;
   wire n_5_2766;
   wire n_5_2767;
   wire n_5_2768;
   wire n_5_2769;
   wire n_5_2770;
   wire n_5_2771;
   wire n_5_2772;
   wire n_5_2773;
   wire n_5_2774;
   wire n_5_2775;
   wire n_5_2776;
   wire n_5_2777;
   wire n_5_2778;
   wire n_5_2779;
   wire n_5_2780;
   wire n_5_2781;
   wire n_5_2782;
   wire n_5_2783;
   wire n_5_2784;
   wire n_5_2785;
   wire n_5_2786;
   wire n_5_2787;
   wire n_5_2788;
   wire n_5_2789;
   wire n_5_2790;
   wire n_5_2791;
   wire n_5_2792;
   wire n_5_2793;
   wire n_5_2794;
   wire n_5_2795;
   wire n_5_2796;
   wire n_5_2797;
   wire n_5_2798;
   wire n_5_2799;
   wire n_5_2800;
   wire n_5_2801;
   wire n_5_2802;
   wire n_5_2803;
   wire n_5_2804;
   wire n_5_2805;
   wire n_5_2806;
   wire n_5_2807;
   wire n_5_2808;
   wire n_5_2809;
   wire n_5_2810;
   wire n_5_2811;
   wire n_5_2812;
   wire n_5_2813;
   wire n_5_2814;
   wire n_5_2815;
   wire n_5_2816;
   wire n_5_2817;
   wire n_5_2818;
   wire n_5_4078;
   wire n_5_2819;
   wire n_5_2820;
   wire n_5_2821;
   wire n_5_2822;
   wire n_5_2823;
   wire n_5_2824;
   wire n_5_2825;
   wire n_5_2826;
   wire n_5_2827;
   wire n_5_2828;
   wire n_5_2829;
   wire n_5_2830;
   wire n_5_2831;
   wire n_5_2832;
   wire n_5_2833;
   wire n_5_2834;
   wire n_5_2835;
   wire n_5_2836;
   wire n_5_2837;
   wire n_5_2838;
   wire n_5_2839;
   wire n_5_2840;
   wire n_5_2841;
   wire n_5_2842;
   wire n_5_2843;
   wire n_5_2844;
   wire n_5_4079;
   wire n_5_2845;
   wire n_5_2846;
   wire n_5_2847;
   wire n_5_2848;
   wire n_5_2849;
   wire n_5_2850;
   wire n_5_2851;
   wire n_5_2852;
   wire n_5_2853;
   wire n_5_2854;
   wire n_5_2855;
   wire n_5_2856;
   wire n_5_2857;
   wire n_5_2858;
   wire n_5_2859;
   wire n_5_2860;
   wire n_5_2861;
   wire n_5_2862;
   wire n_5_2863;
   wire n_5_2864;
   wire n_5_2865;
   wire n_5_2866;
   wire n_5_2867;
   wire n_5_2868;
   wire n_5_2869;
   wire n_5_2870;
   wire n_5_2871;
   wire n_5_2872;
   wire n_5_2873;
   wire n_5_2874;
   wire n_5_2875;
   wire n_5_2876;
   wire n_5_2877;
   wire n_5_2878;
   wire n_5_2879;
   wire n_5_2880;
   wire n_5_2881;
   wire n_5_2882;
   wire n_5_2883;
   wire n_5_2884;
   wire n_5_2885;
   wire n_5_2886;
   wire n_5_2887;
   wire n_5_2888;
   wire n_5_2889;
   wire n_5_2890;
   wire n_5_2891;
   wire n_5_2892;
   wire n_5_2893;
   wire n_5_2894;
   wire n_5_2895;
   wire n_5_2896;
   wire n_5_2897;
   wire n_5_2898;
   wire n_5_2899;
   wire n_5_2900;
   wire n_5_2901;
   wire n_5_2902;
   wire n_5_2903;
   wire n_5_2904;
   wire n_5_2905;
   wire n_5_2906;
   wire n_5_2907;
   wire n_5_2908;
   wire n_5_2909;
   wire n_5_2910;
   wire n_5_2911;
   wire n_5_2912;
   wire n_5_2913;
   wire n_5_2914;
   wire n_5_2915;
   wire n_5_2916;
   wire n_5_2917;
   wire n_5_2918;
   wire n_5_2919;
   wire n_5_2920;
   wire n_5_2921;
   wire n_5_2922;
   wire n_5_2923;
   wire n_5_2924;
   wire n_5_2925;
   wire n_5_4080;
   wire n_5_2926;
   wire n_5_2927;
   wire n_5_4081;
   wire n_5_2928;
   wire n_5_2929;
   wire n_5_2930;
   wire n_5_2931;
   wire n_5_2932;
   wire n_5_2933;
   wire n_5_2934;
   wire n_5_2935;
   wire n_5_2936;
   wire n_5_2937;
   wire n_5_2938;
   wire n_5_2939;
   wire n_5_2940;
   wire n_5_2941;
   wire n_5_2942;
   wire n_5_2943;
   wire n_5_2944;
   wire n_5_2945;
   wire n_5_2946;
   wire n_5_2947;
   wire n_5_2948;
   wire n_5_2949;
   wire n_5_2950;
   wire n_5_2951;
   wire n_5_2952;
   wire n_5_2953;
   wire n_5_2954;
   wire n_5_2955;
   wire n_5_2956;
   wire n_5_2957;
   wire n_5_2958;
   wire n_5_2959;
   wire n_5_2960;
   wire n_5_2961;
   wire n_5_2962;
   wire n_5_2963;
   wire n_5_2964;
   wire n_5_2965;
   wire n_5_3188;
   wire n_5_2966;
   wire n_5_3189;
   wire n_5_2967;
   wire n_5_2968;
   wire n_5_2969;
   wire n_5_2970;
   wire n_5_2971;
   wire n_5_2972;
   wire n_5_2973;
   wire n_5_2974;
   wire n_5_2975;
   wire n_5_2976;
   wire n_5_2977;
   wire n_5_2978;
   wire n_5_2979;
   wire n_5_2980;
   wire n_5_2981;
   wire n_5_2982;
   wire n_5_2983;
   wire n_5_2984;
   wire n_5_2985;
   wire n_5_2986;
   wire n_5_2987;
   wire n_5_2988;
   wire n_5_2989;
   wire n_5_2990;
   wire n_5_2991;
   wire n_5_2992;
   wire n_5_2993;
   wire n_5_2994;
   wire n_5_2995;
   wire n_5_2996;
   wire n_5_2997;
   wire n_5_2998;
   wire n_5_2999;
   wire n_5_3000;
   wire n_5_3001;
   wire n_5_3002;
   wire n_5_3003;
   wire n_5_3004;
   wire n_5_3005;
   wire n_5_3006;
   wire n_5_3007;
   wire n_5_3008;
   wire n_5_3009;
   wire n_5_3010;
   wire n_5_3011;
   wire n_5_3012;
   wire n_5_3013;
   wire n_5_3014;
   wire n_5_3015;
   wire n_5_3016;
   wire n_5_3190;
   wire n_5_3017;
   wire n_5_3018;
   wire n_5_3019;
   wire n_5_3020;
   wire n_5_3021;
   wire n_5_3022;
   wire n_5_3023;
   wire n_5_3024;
   wire n_5_3025;
   wire n_5_3026;
   wire n_5_3027;
   wire n_5_3028;
   wire n_5_3029;
   wire n_5_3030;
   wire n_5_3031;
   wire n_5_3032;
   wire n_5_3033;
   wire n_5_3034;
   wire n_5_3035;
   wire n_5_3036;
   wire n_5_3037;
   wire n_5_3038;
   wire n_5_3039;
   wire n_5_3040;
   wire n_5_3041;
   wire n_5_3042;
   wire n_5_3337;
   wire n_5_3043;
   wire n_5_3044;
   wire n_5_3045;
   wire n_5_3046;
   wire n_5_3047;
   wire n_5_3048;
   wire n_5_3049;
   wire n_5_3050;
   wire n_5_3051;
   wire n_5_3052;
   wire n_5_3053;
   wire n_5_3054;
   wire n_5_3055;
   wire n_5_3056;
   wire n_5_3057;
   wire n_5_3058;
   wire n_5_3059;
   wire n_5_3060;
   wire n_5_3061;
   wire n_5_3062;
   wire n_5_3063;
   wire n_5_3064;
   wire n_5_3065;
   wire n_5_3066;
   wire n_5_3067;
   wire n_5_3068;
   wire n_5_3069;
   wire n_5_3397;
   wire n_5_3070;
   wire n_5_3071;
   wire n_5_3072;
   wire n_5_3073;
   wire n_5_3074;
   wire n_5_3075;
   wire n_5_3076;
   wire n_5_3398;
   wire n_5_3077;
   wire n_5_3078;
   wire n_5_3079;
   wire n_5_3399;
   wire n_5_3080;
   wire n_5_3081;
   wire n_5_3082;
   wire n_5_3083;
   wire n_5_3084;
   wire n_5_3085;
   wire n_5_3086;
   wire n_5_3087;
   wire n_5_3088;
   wire n_5_3089;
   wire n_5_3090;
   wire n_5_3091;
   wire n_5_3092;
   wire n_5_3093;
   wire n_5_3094;
   wire n_5_3095;
   wire n_5_3096;
   wire n_5_3097;
   wire n_5_3098;
   wire n_5_3099;
   wire n_5_3191;
   wire n_5_3100;
   wire n_5_3101;
   wire n_5_3102;
   wire n_5_3103;
   wire n_5_3104;
   wire n_5_3105;
   wire n_5_3106;
   wire n_5_3107;
   wire n_5_3108;
   wire n_5_3109;
   wire n_5_3110;
   wire n_5_3111;
   wire n_5_3112;
   wire n_5_3113;
   wire n_5_3114;
   wire n_5_3115;
   wire n_5_3116;
   wire n_5_3117;
   wire n_5_3118;
   wire n_5_3119;
   wire n_5_3120;
   wire n_5_3121;
   wire n_5_3122;
   wire n_5_3123;
   wire n_5_3125;
   wire n_5_3127;
   wire n_5_3130;
   wire n_5_3132;
   wire n_5_3133;
   wire n_5_3134;
   wire n_5_3135;
   wire n_5_3137;
   wire n_5_3140;
   wire n_5_3144;
   wire n_5_3145;
   wire n_5_3146;
   wire n_5_3150;
   wire n_5_3153;
   wire n_5_3154;
   wire n_5_3155;
   wire n_5_3156;
   wire n_5_3159;
   wire n_5_3161;
   wire n_5_3169;
   wire n_5_3184;
   wire n_5_3186;
   wire n_5_3187;
   wire n_5_3192;
   wire n_5_3193;
   wire n_5_3194;
   wire n_5_3195;
   wire n_5_3196;
   wire n_5_3197;
   wire n_5_3198;
   wire n_5_4082;
   wire n_5_4083;
   wire n_5_4084;
   wire n_5_3199;
   wire n_5_3200;
   wire n_5_3201;
   wire n_5_3202;
   wire n_5_3203;
   wire n_5_3204;
   wire n_5_3205;
   wire n_5_3206;
   wire n_5_3207;
   wire n_5_3208;
   wire n_5_3209;
   wire n_5_3210;
   wire n_5_3211;
   wire n_5_3212;
   wire n_5_3213;
   wire n_5_3214;
   wire n_5_3215;
   wire n_5_3216;
   wire n_5_3217;
   wire n_5_3218;
   wire n_5_3219;
   wire n_5_3220;
   wire n_5_3221;
   wire n_5_3222;
   wire n_5_3223;
   wire n_5_3224;
   wire n_5_3225;
   wire n_5_3226;
   wire n_5_3227;
   wire n_5_3228;
   wire n_5_3229;
   wire n_5_3230;
   wire n_5_3231;
   wire n_5_3232;
   wire n_5_3233;
   wire n_5_3234;
   wire n_5_3235;
   wire n_5_3236;
   wire n_5_3237;
   wire n_5_3238;
   wire n_5_3239;
   wire n_5_3240;
   wire n_5_3241;
   wire n_5_3242;
   wire n_5_3243;
   wire n_5_3244;
   wire n_5_3245;
   wire n_5_3246;
   wire n_5_3247;
   wire n_5_3248;
   wire n_5_3249;
   wire n_5_4085;
   wire n_5_3250;
   wire n_5_3251;
   wire n_5_3252;
   wire n_5_3253;
   wire n_5_3254;
   wire n_5_3255;
   wire n_5_3256;
   wire n_5_3257;
   wire n_5_3258;
   wire n_5_3259;
   wire n_5_3260;
   wire n_5_3261;
   wire n_5_3262;
   wire n_5_3263;
   wire n_5_3264;
   wire n_5_3265;
   wire n_5_3266;
   wire n_5_3267;
   wire n_5_3268;
   wire n_5_3269;
   wire n_5_3270;
   wire n_5_3271;
   wire n_5_3272;
   wire n_5_3273;
   wire n_5_3274;
   wire n_5_3275;
   wire n_5_3276;
   wire n_5_3277;
   wire n_5_3278;
   wire n_5_3279;
   wire n_5_3280;
   wire n_5_3281;
   wire n_5_3282;
   wire n_5_3283;
   wire n_5_3284;
   wire n_5_3285;
   wire n_5_3286;
   wire n_5_3287;
   wire n_5_3288;
   wire n_5_3289;
   wire n_5_3290;
   wire n_5_3291;
   wire n_5_3292;
   wire n_5_3293;
   wire n_5_3294;
   wire n_5_3295;
   wire n_5_3296;
   wire n_5_3297;
   wire n_5_3298;
   wire n_5_3299;
   wire n_5_3300;
   wire n_5_3301;
   wire n_5_3302;
   wire n_5_3303;
   wire n_5_3304;
   wire n_5_3305;
   wire n_5_3306;
   wire n_5_3307;
   wire n_5_3308;
   wire n_5_3309;
   wire n_5_3310;
   wire n_5_3311;
   wire n_5_3312;
   wire n_5_3313;
   wire n_5_3314;
   wire n_5_3315;
   wire n_5_3316;
   wire n_5_3401;
   wire n_5_3317;
   wire n_5_3318;
   wire n_5_3319;
   wire n_5_3320;
   wire n_5_3321;
   wire n_5_3322;
   wire n_5_3323;
   wire n_5_3324;
   wire n_5_3325;
   wire n_5_3326;
   wire n_5_3327;
   wire n_5_3328;
   wire n_5_3329;
   wire n_5_3330;
   wire n_5_3331;
   wire n_5_3334;
   wire n_5_3336;
   wire n_5_3342;
   wire n_5_3344;
   wire n_5_3346;
   wire n_5_3348;
   wire n_5_3349;
   wire n_5_3351;
   wire n_5_3403;
   wire n_5_462;
   wire n_5_3354;
   wire n_5_3358;
   wire n_5_3361;
   wire n_5_3362;
   wire n_5_3363;
   wire n_5_3368;
   wire n_5_3369;
   wire n_5_3370;
   wire n_5_3371;
   wire n_5_3373;
   wire n_5_3374;
   wire n_5_3375;
   wire n_5_3376;
   wire n_5_3378;
   wire n_5_3382;
   wire n_5_3388;
   wire n_5_3390;
   wire n_5_3391;
   wire n_5_3394;
   wire n_5_3395;
   wire n_5_3396;
   wire n_5_3400;
   wire n_5_3402;
   wire n_5_3404;
   wire n_5_3405;
   wire n_5_3406;
   wire n_5_3407;
   wire n_5_3408;
   wire n_5_3409;
   wire n_5_3410;
   wire n_5_3411;
   wire n_5_3412;
   wire n_5_3413;
   wire n_5_3414;
   wire n_5_3415;
   wire n_5_3416;
   wire n_5_3417;
   wire n_5_3418;
   wire n_5_3419;
   wire n_5_3420;
   wire n_5_3421;
   wire n_5_3422;
   wire n_5_3423;
   wire n_5_3424;
   wire n_5_3425;
   wire n_5_3426;
   wire n_5_3427;
   wire n_5_3428;
   wire n_5_3429;
   wire n_5_3430;
   wire n_5_3431;
   wire n_5_3432;
   wire n_5_3433;
   wire n_5_3434;
   wire n_5_3435;
   wire n_5_3436;
   wire n_5_3437;
   wire n_5_3438;
   wire n_5_3439;
   wire n_5_3440;
   wire n_5_3441;
   wire n_5_3442;
   wire n_5_4086;
   wire n_5_4087;
   wire n_5_3443;
   wire n_5_3444;
   wire n_5_3445;
   wire n_5_3446;
   wire n_5_3447;
   wire n_5_3448;
   wire n_5_3449;
   wire n_5_3450;
   wire n_5_3451;
   wire n_5_3452;
   wire n_5_3453;
   wire n_5_3454;
   wire n_5_3455;
   wire n_5_3456;
   wire n_5_3457;
   wire n_5_3458;
   wire n_5_3459;
   wire n_5_3460;
   wire n_5_3461;
   wire n_5_3462;
   wire n_5_3463;
   wire n_5_3464;
   wire n_5_3465;
   wire n_5_3466;
   wire n_5_3467;
   wire n_5_3468;
   wire n_5_3469;
   wire n_5_3470;
   wire n_5_3471;
   wire n_5_3472;
   wire n_5_3473;
   wire n_5_3474;
   wire n_5_3475;
   wire n_5_3476;
   wire n_5_3477;
   wire n_5_3478;
   wire n_5_3479;
   wire n_5_3480;
   wire n_5_3481;
   wire n_5_3482;
   wire n_5_3483;
   wire n_5_3484;
   wire n_5_3485;
   wire n_5_3486;
   wire n_5_3487;
   wire n_5_3488;
   wire n_5_3489;
   wire n_5_3490;
   wire n_5_3491;
   wire n_5_3492;
   wire n_5_3493;
   wire n_5_3494;
   wire n_5_3495;
   wire n_5_3496;
   wire n_5_3497;
   wire n_5_3498;
   wire n_5_3499;
   wire n_5_4088;
   wire n_5_3500;
   wire n_5_3501;
   wire n_5_3502;
   wire n_5_3503;
   wire n_5_3504;
   wire n_5_3505;
   wire n_5_3506;
   wire n_5_3507;
   wire n_5_3508;
   wire n_5_3509;
   wire n_5_3510;
   wire n_5_3511;
   wire n_5_3512;
   wire n_5_3513;
   wire n_5_3514;
   wire n_5_3515;
   wire n_5_3516;
   wire n_5_3517;
   wire n_5_3518;
   wire n_5_3519;
   wire n_5_3520;
   wire n_5_3521;
   wire n_5_3522;
   wire n_5_3523;
   wire n_5_3524;
   wire n_5_3525;
   wire n_5_3526;
   wire n_5_3527;
   wire n_5_3528;
   wire n_5_3529;
   wire n_5_3530;
   wire n_5_464;
   wire n_5_3532;
   wire n_5_3533;
   wire n_5_3534;
   wire n_5_3535;
   wire n_5_3536;
   wire n_5_3537;
   wire n_5_3538;
   wire n_5_3539;
   wire n_5_3540;
   wire n_5_3541;
   wire n_5_3542;
   wire n_5_3543;
   wire n_5_3544;
   wire n_5_3545;
   wire n_5_3546;
   wire n_5_3547;
   wire n_5_3548;
   wire n_5_3549;
   wire n_5_3550;
   wire n_5_3551;
   wire n_5_3552;
   wire n_5_3553;
   wire n_5_3554;
   wire n_5_3555;
   wire n_5_3556;
   wire n_5_3557;
   wire n_5_3558;
   wire n_5_3559;
   wire n_5_3560;
   wire n_5_3561;
   wire n_5_3562;
   wire n_5_3563;
   wire n_5_3564;
   wire n_5_3565;
   wire n_5_3566;
   wire n_5_3567;
   wire n_5_4656;
   wire n_5_4657;
   wire n_5_3568;
   wire n_5_3569;
   wire n_5_3570;
   wire n_5_3571;
   wire n_5_3572;
   wire n_5_3573;
   wire n_5_3574;
   wire n_5_3575;
   wire n_5_3576;
   wire n_5_3577;
   wire n_5_3578;
   wire n_5_3579;
   wire n_5_3580;
   wire n_5_3581;
   wire n_5_3582;
   wire n_5_3583;
   wire n_5_3584;
   wire n_5_3585;
   wire n_5_3586;
   wire n_5_4089;
   wire n_5_3587;
   wire n_5_4090;
   wire n_5_3588;
   wire n_5_4091;
   wire n_5_3589;
   wire n_5_4092;
   wire n_5_4093;
   wire n_5_3590;
   wire n_5_3591;
   wire n_5_3592;
   wire n_5_3593;
   wire n_5_3594;
   wire n_5_3595;
   wire n_5_3596;
   wire n_5_3597;
   wire n_5_3598;
   wire n_5_3599;
   wire n_5_3600;
   wire n_5_3601;
   wire n_5_3602;
   wire n_5_3603;
   wire n_5_4094;
   wire n_5_3604;
   wire n_5_3605;
   wire n_5_3606;
   wire n_5_3607;
   wire n_5_3608;
   wire n_5_3609;
   wire n_5_3610;
   wire n_5_3611;
   wire n_5_3612;
   wire n_5_3613;
   wire n_5_3614;
   wire n_5_3615;
   wire n_5_3616;
   wire n_5_3617;
   wire n_5_3618;
   wire n_5_3619;
   wire n_5_3620;
   wire n_5_3621;
   wire n_5_3622;
   wire n_5_3623;
   wire n_5_3624;
   wire n_5_4095;
   wire n_5_3625;
   wire n_5_3626;
   wire n_5_3627;
   wire n_5_3628;
   wire n_5_3629;
   wire n_5_3630;
   wire n_5_3631;
   wire n_5_3633;
   wire n_5_4096;
   wire n_5_3634;
   wire n_5_3635;
   wire n_5_3636;
   wire n_5_3637;
   wire n_5_3638;
   wire n_5_3640;
   wire n_5_3641;
   wire n_5_3642;
   wire n_5_3643;
   wire n_5_3644;
   wire n_5_3645;
   wire n_5_3646;
   wire n_5_3647;
   wire n_5_3648;
   wire n_5_3649;
   wire n_5_3650;
   wire n_5_3651;
   wire n_5_3652;
   wire n_5_3653;
   wire n_5_3654;
   wire n_5_3655;
   wire n_5_4097;
   wire n_5_3656;
   wire n_5_3657;
   wire n_5_3658;
   wire n_5_3659;
   wire n_5_3660;
   wire n_5_3661;
   wire n_5_3662;
   wire n_5_3663;
   wire n_5_3664;
   wire n_5_4098;
   wire n_5_3665;
   wire n_5_3666;
   wire n_5_3667;
   wire n_5_3668;
   wire n_5_3669;
   wire n_5_3670;
   wire n_5_3671;
   wire n_5_3672;
   wire n_5_3673;
   wire n_5_3674;
   wire n_5_3675;
   wire n_5_3676;
   wire n_5_3677;
   wire n_5_3678;
   wire n_5_3679;
   wire n_5_4099;
   wire n_5_3680;
   wire n_5_3683;
   wire n_5_3684;
   wire n_5_3685;
   wire n_5_3686;
   wire n_5_3687;
   wire n_5_3688;
   wire n_5_3689;
   wire n_5_3690;
   wire n_5_3691;
   wire n_5_3692;
   wire n_5_3693;
   wire n_5_3694;
   wire n_5_3695;
   wire n_5_3696;
   wire n_5_3697;
   wire n_5_3698;
   wire n_5_3699;
   wire n_5_3700;
   wire n_5_3701;
   wire n_5_3702;
   wire n_5_3703;
   wire n_5_3704;
   wire n_5_476;
   wire n_5_486;
   wire n_5_497;
   wire n_5_4100;
   wire n_5_3711;
   wire n_5_3712;
   wire n_5_3713;
   wire n_5_3714;
   wire n_5_3715;
   wire n_5_3716;
   wire n_5_3717;
   wire n_5_3718;
   wire n_5_3719;
   wire n_5_3720;
   wire n_5_3721;
   wire n_5_3722;
   wire n_5_3723;
   wire n_5_3724;
   wire n_5_3725;
   wire n_5_3726;
   wire n_5_3727;
   wire n_5_3728;
   wire n_5_3729;
   wire n_5_3730;
   wire n_5_3731;
   wire n_5_3732;
   wire n_5_3733;
   wire n_5_3734;
   wire n_5_3735;
   wire n_5_3737;
   wire n_5_3738;
   wire n_5_3739;
   wire n_5_3740;
   wire n_5_3741;
   wire n_5_3742;
   wire n_5_3743;
   wire n_5_3744;
   wire n_5_3745;
   wire n_5_3746;
   wire n_5_3747;
   wire n_5_4658;
   wire n_5_3748;
   wire n_5_3749;
   wire n_5_3750;
   wire n_5_3751;
   wire n_5_4101;
   wire n_5_3752;
   wire n_5_4659;
   wire n_5_3753;
   wire n_5_3754;
   wire n_5_3755;
   wire n_5_4102;
   wire n_5_3756;
   wire n_5_3757;
   wire n_5_3758;
   wire n_5_4103;
   wire n_5_3759;
   wire n_5_3760;
   wire n_5_3761;
   wire n_5_3762;
   wire n_5_3763;
   wire n_5_3764;
   wire n_5_3765;
   wire n_5_3766;
   wire n_5_3767;
   wire n_5_3768;
   wire n_5_3769;
   wire n_5_3770;
   wire n_5_873;
   wire n_5_3772;
   wire n_5_3773;
   wire n_5_3774;
   wire n_5_3775;
   wire n_5_3776;
   wire n_5_3777;
   wire n_5_3778;
   wire n_5_4104;
   wire n_5_3779;
   wire n_5_3780;
   wire n_5_3781;
   wire n_5_3782;
   wire n_5_3783;
   wire n_5_3784;
   wire n_5_3785;
   wire n_5_3786;
   wire n_5_3787;
   wire n_5_3788;
   wire n_5_3789;
   wire n_5_3790;
   wire n_5_3791;
   wire n_5_3792;
   wire n_5_3793;
   wire n_5_3794;
   wire n_5_3795;
   wire n_5_3796;
   wire n_5_3797;
   wire n_5_3798;
   wire n_5_3799;
   wire n_5_3865;
   wire n_5_3800;
   wire n_5_3801;
   wire n_5_3802;
   wire n_5_3803;
   wire n_5_3804;
   wire n_5_3805;
   wire n_5_498;
   wire n_5_3810;
   wire n_5_3811;
   wire n_5_3812;
   wire n_5_3813;
   wire n_5_3814;
   wire n_5_3815;
   wire n_5_3816;
   wire n_5_3817;
   wire n_5_3818;
   wire n_5_3819;
   wire n_5_3820;
   wire n_5_3821;
   wire n_5_3822;
   wire n_5_3823;
   wire n_5_3824;
   wire n_5_3825;
   wire n_5_3826;
   wire n_5_4107;
   wire n_5_3827;
   wire n_5_3828;
   wire n_5_3829;
   wire n_5_3830;
   wire n_5_3831;
   wire n_5_3832;
   wire n_5_3833;
   wire n_5_3834;
   wire n_5_3835;
   wire n_5_3836;
   wire n_5_3837;
   wire n_5_3838;
   wire n_5_3842;
   wire n_5_3843;
   wire n_5_3844;
   wire n_5_3845;
   wire n_5_3846;
   wire n_5_3847;
   wire n_5_3848;
   wire n_5_3849;
   wire n_5_3850;
   wire n_5_4108;
   wire n_5_3851;
   wire n_5_3852;
   wire n_5_3853;
   wire n_5_3854;
   wire n_5_3870;
   wire n_5_3884;
   wire n_5_3885;
   wire n_5_3892;
   wire n_5_3894;
   wire n_5_3896;
   wire n_5_3900;
   wire n_5_3901;
   wire n_5_3902;
   wire n_5_4109;
   wire n_5_3908;
   wire n_5_3909;
   wire n_5_3915;
   wire n_5_3917;
   wire n_5_3919;
   wire n_5_3924;
   wire n_5_3926;
   wire n_5_3929;
   wire n_5_3933;
   wire n_5_3958;
   wire n_5_3962;
   wire n_5_3980;
   wire n_5_3981;
   wire n_5_3986;
   wire n_5_3988;
   wire n_5_3992;
   wire n_5_4000;
   wire n_5_4004;
   wire n_5_4014;
   wire n_5_4110;
   wire n_5_4111;
   wire n_5_4018;
   wire n_5_4046;
   wire n_5_4047;
   wire n_5_4112;
   wire n_5_4054;
   wire n_5_4105;
   wire n_5_4106;
   wire n_5_4113;
   wire n_5_4114;
   wire n_5_4115;
   wire n_5_4116;
   wire n_5_4117;
   wire n_5_4118;
   wire n_5_4119;
   wire n_5_4120;
   wire n_5_4121;
   wire n_5_4122;
   wire n_5_4123;
   wire n_5_4124;
   wire n_5_4125;
   wire n_5_4126;
   wire n_5_4127;
   wire n_5_4128;
   wire n_5_4129;
   wire n_5_4130;
   wire n_5_4131;
   wire n_5_4132;
   wire n_5_4133;
   wire n_5_4134;
   wire n_5_4135;
   wire n_5_4136;
   wire n_5_4137;
   wire n_5_4138;
   wire n_5_4139;
   wire n_5_4140;
   wire n_5_515;
   wire n_5_4141;
   wire n_5_4142;
   wire n_5_4143;
   wire n_5_4144;
   wire n_5_4145;
   wire n_5_4146;
   wire n_5_4147;
   wire n_5_4148;
   wire n_5_4149;
   wire n_5_4150;
   wire n_5_4151;
   wire n_5_4152;
   wire n_5_4153;
   wire n_5_4154;
   wire n_5_4155;
   wire n_5_4156;
   wire n_5_4157;
   wire n_5_4158;
   wire n_5_4159;
   wire n_5_4160;
   wire n_5_4161;
   wire n_5_4162;
   wire n_5_4163;
   wire n_5_4164;
   wire n_5_4165;
   wire n_5_4166;
   wire n_5_4167;
   wire n_5_4168;
   wire n_5_4169;
   wire n_5_4170;
   wire n_5_4171;
   wire n_5_4172;
   wire n_5_4173;
   wire n_5_4174;
   wire n_5_4175;
   wire n_5_4176;
   wire n_5_4177;
   wire n_5_4178;
   wire n_5_4179;
   wire n_5_4180;
   wire n_5_4181;
   wire n_5_4182;
   wire n_5_4183;
   wire n_5_4184;
   wire n_5_4185;
   wire n_5_4186;
   wire n_5_4187;
   wire n_5_4188;
   wire n_5_4189;
   wire n_5_4190;
   wire n_5_4191;
   wire n_5_4192;
   wire n_5_4193;
   wire n_5_4194;
   wire n_5_4195;
   wire n_5_4196;
   wire n_5_4197;
   wire n_5_4198;
   wire n_5_4199;
   wire n_5_4200;
   wire n_5_4201;
   wire n_5_4202;
   wire n_5_4203;
   wire n_5_4204;
   wire n_5_4205;
   wire n_5_4206;
   wire n_5_4207;
   wire n_5_4208;
   wire n_5_4209;
   wire n_5_4210;
   wire n_5_4211;
   wire n_5_4212;
   wire n_5_4213;
   wire n_5_4214;
   wire n_5_4215;
   wire n_5_4216;
   wire n_5_4217;
   wire n_5_4218;
   wire n_5_4219;
   wire n_5_4220;
   wire n_5_4221;
   wire n_5_524;
   wire n_5_4223;
   wire n_5_4663;
   wire n_5_4224;
   wire n_5_4225;
   wire n_5_4226;
   wire n_5_4227;
   wire n_5_4228;
   wire n_5_4229;
   wire n_5_4230;
   wire n_5_525;
   wire n_5_4232;
   wire n_5_4233;
   wire n_5_4234;
   wire n_5_4235;
   wire n_5_4236;
   wire n_5_4237;
   wire n_5_4238;
   wire n_5_4239;
   wire n_5_4240;
   wire n_5_4241;
   wire n_5_4242;
   wire n_5_526;
   wire n_5_4243;
   wire n_5_4244;
   wire n_5_4245;
   wire n_5_4246;
   wire n_5_4248;
   wire n_5_4249;
   wire n_5_4250;
   wire n_5_4251;
   wire n_5_4252;
   wire n_5_4253;
   wire n_5_4254;
   wire n_5_4256;
   wire n_5_4257;
   wire n_5_528;
   wire n_5_576;
   wire n_5_622;
   wire n_5_4262;
   wire n_5_4263;
   wire n_5_4264;
   wire n_5_4265;
   wire n_5_4266;
   wire n_5_531;
   wire n_5_4269;
   wire n_5_4270;
   wire n_5_4271;
   wire n_5_4272;
   wire n_5_4273;
   wire n_5_4274;
   wire n_5_4275;
   wire n_5_4276;
   wire n_5_4277;
   wire n_5_4278;
   wire n_5_4280;
   wire n_5_4281;
   wire n_5_4282;
   wire n_5_4283;
   wire n_5_4284;
   wire n_5_4285;
   wire n_5_4286;
   wire n_5_4287;
   wire n_5_4288;
   wire n_5_4289;
   wire n_5_4290;
   wire n_5_4292;
   wire n_5_4293;
   wire n_5_4294;
   wire n_5_4295;
   wire n_5_4296;
   wire n_5_4297;
   wire n_5_532;
   wire n_5_4299;
   wire n_5_4300;
   wire n_5_536;
   wire n_5_4302;
   wire n_5_4303;
   wire n_5_4304;
   wire n_5_4305;
   wire n_5_4306;
   wire n_5_215;
   wire n_5_4308;
   wire n_5_4309;
   wire n_5_216;
   wire n_5_4311;
   wire n_5_4312;
   wire n_5_4313;
   wire n_5_4314;
   wire n_5_4315;
   wire n_5_4316;
   wire n_5_4317;
   wire n_5_4318;
   wire n_5_4319;
   wire n_5_3873;
   wire n_5_4321;
   wire n_5_4322;
   wire n_5_4323;
   wire n_5_4324;
   wire n_5_4325;
   wire n_5_4329;
   wire n_5_4330;
   wire n_5_4331;
   wire n_5_4332;
   wire n_5_4333;
   wire n_5_4334;
   wire n_5_4335;
   wire n_5_4336;
   wire n_5_4337;
   wire n_5_4338;
   wire n_5_4339;
   wire n_5_4340;
   wire n_5_4341;
   wire n_5_4342;
   wire n_5_4343;
   wire n_5_4346;
   wire n_5_4347;
   wire n_5_4348;
   wire n_5_219;
   wire n_5_4350;
   wire n_5_4351;
   wire n_5_4352;
   wire n_5_4353;
   wire n_5_539;
   wire n_5_4355;
   wire n_5_4356;
   wire n_5_4357;
   wire n_5_4358;
   wire n_5_4359;
   wire n_5_4360;
   wire n_5_4361;
   wire n_5_4364;
   wire n_5_4365;
   wire n_5_4366;
   wire n_5_4367;
   wire n_5_4368;
   wire n_5_546;
   wire n_5_578;
   wire n_5_4373;
   wire n_5_4374;
   wire n_5_4375;
   wire n_5_4376;
   wire n_5_4377;
   wire n_5_4378;
   wire n_5_4379;
   wire n_5_579;
   wire n_5_581;
   wire n_5_4383;
   wire n_5_4384;
   wire n_5_4385;
   wire n_5_4386;
   wire n_5_4387;
   wire n_5_4388;
   wire n_5_4389;
   wire n_5_4392;
   wire n_5_4393;
   wire n_5_4394;
   wire n_5_4395;
   wire n_5_4396;
   wire n_5_4397;
   wire n_5_4398;
   wire n_5_4399;
   wire n_5_4400;
   wire n_5_4401;
   wire n_5_4402;
   wire n_5_4403;
   wire n_5_4404;
   wire n_5_616;
   wire n_5_4406;
   wire n_5_4407;
   wire n_5_4408;
   wire n_5_625;
   wire n_5_4412;
   wire n_5_4413;
   wire n_5_4414;
   wire n_5_4415;
   wire n_5_4416;
   wire n_5_4417;
   wire n_5_626;
   wire n_5_646;
   wire n_5_4422;
   wire n_5_4423;
   wire n_5_4424;
   wire n_5_4425;
   wire n_5_4426;
   wire n_5_4427;
   wire n_5_4428;
   wire n_5_4429;
   wire n_5_4430;
   wire n_5_4431;
   wire n_5_4432;
   wire n_5_4433;
   wire n_5_4434;
   wire n_5_4435;
   wire n_5_4436;
   wire n_5_4437;
   wire n_5_4438;
   wire n_5_647;
   wire n_5_4440;
   wire n_5_4441;
   wire n_5_4442;
   wire n_5_4443;
   wire n_5_4444;
   wire n_5_4445;
   wire n_5_4446;
   wire n_5_876;
   wire n_5_4448;
   wire n_5_4449;
   wire n_5_4450;
   wire n_5_4451;
   wire n_5_4452;
   wire n_5_4453;
   wire n_5_4454;
   wire n_5_4455;
   wire n_5_4456;
   wire n_5_4457;
   wire n_5_4458;
   wire n_5_256;
   wire n_5_4460;
   wire n_5_4461;
   wire n_5_4462;
   wire n_5_4463;
   wire n_5_4464;
   wire n_5_4465;
   wire n_5_4466;
   wire n_5_4467;
   wire n_5_4468;
   wire n_5_4469;
   wire n_5_4470;
   wire n_5_4471;
   wire n_5_4472;
   wire n_5_4473;
   wire n_5_4474;
   wire n_5_4475;
   wire n_5_4476;
   wire n_5_4477;
   wire n_5_4478;
   wire n_5_4479;
   wire n_5_4480;
   wire n_5_4481;
   wire n_5_4482;
   wire n_5_4483;
   wire n_5_4484;
   wire n_5_4486;
   wire n_5_4487;
   wire n_5_4488;
   wire n_5_4489;
   wire n_5_4490;
   wire n_5_4670;
   wire n_5_4492;
   wire n_5_4493;
   wire n_5_4495;
   wire n_5_4496;
   wire n_5_4497;
   wire n_5_4498;
   wire n_5_4499;
   wire n_5_4500;
   wire n_5_4501;
   wire n_5_294;
   wire n_5_4503;
   wire n_5_4504;
   wire n_5_4505;
   wire n_5_4506;
   wire n_5_4507;
   wire n_5_4508;
   wire n_5_649;
   wire n_5_4510;
   wire n_5_4511;
   wire n_5_4512;
   wire n_5_4513;
   wire n_5_4514;
   wire n_5_4515;
   wire n_5_4516;
   wire n_5_4517;
   wire n_5_4518;
   wire n_5_4519;
   wire n_5_4520;
   wire n_5_291;
   wire n_5_4522;
   wire n_5_316;
   wire n_5_4524;
   wire n_5_4526;
   wire n_5_4527;
   wire n_5_4528;
   wire n_5_4529;
   wire n_5_4530;
   wire n_5_4531;
   wire n_5_678;
   wire n_5_4533;
   wire n_5_4534;
   wire n_5_4538;
   wire n_5_4671;
   wire n_5_684;
   wire n_5_692;
   wire n_5_3890;
   wire n_5_4548;
   wire n_5_4549;
   wire n_5_4553;
   wire n_5_4554;
   wire n_5_4672;
   wire n_5_4559;
   wire n_5_4560;
   wire n_5_4561;
   wire n_5_4562;
   wire n_5_4563;
   wire n_5_4564;
   wire n_5_4565;
   wire n_5_4566;
   wire n_5_432;
   wire n_5_4568;
   wire n_5_4569;
   wire n_5_4570;
   wire n_5_443;
   wire n_5_4573;
   wire n_5_4574;
   wire n_5_4575;
   wire n_5_700;
   wire n_5_4577;
   wire n_5_4673;
   wire n_5_429;
   wire n_5_4580;
   wire n_5_4581;
   wire n_5_4582;
   wire n_5_4583;
   wire n_5_4584;
   wire n_5_4585;
   wire n_5_4586;
   wire n_5_4587;
   wire n_5_4588;
   wire n_5_4674;
   wire n_5_4675;
   wire n_5_4676;
   wire n_5_4677;
   wire n_5_4678;
   wire n_5_4679;
   wire n_5_4680;
   wire n_5_4681;
   wire n_5_4682;
   wire n_5_4683;
   wire n_5_4684;
   wire n_5_4685;
   wire n_5_4686;
   wire n_5_4687;
   wire n_5_4688;
   wire n_5_4689;
   wire n_5_4690;
   wire n_5_701;
   wire n_5_4694;
   wire n_5_4695;
   wire n_5_4696;
   wire n_5_4697;
   wire n_5_4698;
   wire n_5_4699;
   wire n_5_4700;
   wire n_5_4702;
   wire n_5_4703;
   wire n_5_4704;
   wire n_5_4589;
   wire n_5_4705;
   wire n_5_4706;
   wire n_5_4707;
   wire n_5_4709;
   wire n_5_465;
   wire n_5_4711;
   wire n_5_4712;
   wire n_5_4713;
   wire n_5_4714;
   wire n_5_4715;
   wire n_5_702;
   wire n_5_4718;
   wire n_5_711;
   wire n_5_716;
   wire n_5_728;
   wire n_5_739;
   wire n_5_3705;
   wire n_5_4728;
   wire n_5_4729;
   wire n_5_4730;
   wire n_5_4731;
   wire n_5_4732;
   wire n_5_3706;
   wire n_5_4734;
   wire n_5_3856;
   wire n_5_749;
   wire n_5_821;
   wire n_5_1031;
   wire n_5_1032;
   wire n_5_1373;
   wire n_5_1374;
   wire n_5_1382;
   wire n_5_2184;
   wire n_5_3353;
   wire n_5_3531;
   wire n_5_3632;
   wire n_5_3639;
   wire n_5_3681;
   wire n_5_3707;
   wire n_5_3708;
   wire n_5_3709;
   wire n_5_3710;
   wire n_5_3806;
   wire n_5_3807;
   wire n_5_3809;
   wire n_5_3871;
   wire n_5_3872;
   wire n_5_3874;
   wire n_5_3875;
   wire n_5_3876;
   wire n_5_3878;
   wire n_5_3930;
   wire n_5_3895;
   wire n_5_3897;
   wire n_5_3899;
   wire n_5_3911;
   wire n_5_3912;
   wire n_5_3913;
   wire n_5_3914;
   wire n_5_3922;
   wire n_5_3923;
   wire n_5_3925;
   wire n_5_3945;
   wire n_5_3956;
   wire n_5_3960;
   wire n_5_3983;
   wire n_5_3984;
   wire n_5_3985;
   wire n_5_3857;
   wire n_5_3997;
   wire n_5_4008;
   wire n_5_4009;
   wire n_5_4055;
   wire n_5_4058;
   wire n_5_4231;
   wire n_5_4247;
   wire n_5_4255;
   wire n_5_4258;
   wire n_5_4261;
   wire n_5_4267;
   wire n_5_4268;
   wire n_5_4291;
   wire n_5_4298;
   wire n_5_4301;
   wire n_5_4354;
   wire n_5_4362;
   wire n_5_4363;
   wire n_5_4369;
   wire n_5_4370;
   wire n_5_4371;
   wire n_5_4380;
   wire n_5_4381;
   wire n_5_4382;
   wire n_5_4390;
   wire n_5_4391;
   wire n_5_4405;
   wire n_5_4409;
   wire n_5_4410;
   wire n_5_4411;
   wire n_5_4418;
   wire n_5_4419;
   wire n_5_4420;
   wire n_5_4421;
   wire n_5_4439;
   wire n_5_4485;
   wire n_5_3931;
   wire n_5_4509;
   wire n_5_4532;
   wire n_5_4535;
   wire n_5_4536;
   wire n_5_4537;
   wire n_5_4539;
   wire n_5_3932;
   wire n_5_3935;
   wire n_5_4543;
   wire n_5_3936;
   wire n_5_4551;
   wire n_5_4552;
   wire n_5_3858;
   wire n_5_3961;
   wire n_5_4557;
   wire n_5_4558;
   wire n_5_4576;
   wire n_5_4578;
   wire n_5_4590;
   wire n_5_4597;
   wire n_5_4602;
   wire n_5_3859;
   wire n_5_4609;
   wire n_5_4610;
   wire n_5_4617;
   wire n_5_4618;
   wire n_5_4619;
   wire n_5_4623;
   wire n_5_3860;
   wire n_5_4625;
   wire n_5_4628;
   wire n_5_4629;
   wire n_5_4630;
   wire n_5_4638;
   wire n_5_4643;
   wire n_5_4650;
   wire n_5_4651;
   wire n_5_4652;
   wire n_5_4660;
   wire n_5_4661;
   wire n_5_4662;
   wire n_5_4664;
   wire n_5_4665;
   wire n_5_4666;
   wire n_5_4667;
   wire n_5_4668;
   wire n_5_4691;
   wire n_5_4692;
   wire n_5_4693;
   wire n_5_4708;
   wire n_5_4716;
   wire n_5_4717;
   wire n_5_4719;
   wire n_5_4722;
   wire n_5_4723;
   wire n_5_3861;
   wire n_5_4725;
   wire n_5_4736;
   wire n_5_4737;
   wire n_5_4738;
   wire n_5_4739;
   wire n_5_4740;
   wire n_5_4741;
   wire n_5_4742;
   wire n_5_4743;
   wire n_5_4744;
   wire n_5_4745;
   wire n_5_4746;
   wire n_5_4747;
   wire n_5_4748;
   wire n_5_4749;
   wire n_5_4750;
   wire n_5_4751;
   wire n_5_4752;
   wire n_5_878;
   wire n_5_4754;
   wire n_5_4755;
   wire n_5_4756;
   wire n_5_4757;
   wire n_5_4758;
   wire n_5_4759;
   wire n_5_4760;
   wire n_5_4761;
   wire n_5_4762;
   wire n_5_4763;
   wire n_5_4764;
   wire n_5_4765;
   wire n_5_4766;
   wire n_5_4767;
   wire n_5_4768;
   wire n_5_4259;
   wire n_5_4260;
   wire n_5_4279;
   wire n_5_4320;
   wire n_5_4774;
   wire n_5_4775;
   wire n_5_4776;
   wire n_5_4777;
   wire n_5_4778;
   wire n_5_4779;
   wire n_5_4780;
   wire n_5_4781;
   wire n_5_4782;
   wire n_5_4783;
   wire n_5_4784;
   wire n_5_4785;
   wire n_5_4786;
   wire n_5_4787;
   wire n_5_4788;
   wire n_5_4789;
   wire n_5_619;
   wire n_5_843;
   wire n_5_3937;
   wire n_5_4037;
   wire n_5_4040;
   wire n_5_4525;
   wire n_5_4579;
   wire n_5_4790;
   wire n_5_4791;
   wire n_5_3771;
   wire n_5_3839;
   wire n_5_3840;
   wire n_5_3841;
   wire n_5_3959;
   wire n_5_3982;
   wire n_5_4222;
   wire n_5_4447;
   wire n_5_4600;
   wire n_5_4613;
   wire n_5_4654;
   wire n_5_4701;
   wire n_5_4753;
   wire n_5_4792;
   wire n_5_4793;
   wire n_5_4794;
   wire n_5_4795;
   wire n_5_4326;
   wire n_5_4327;
   wire n_5_4328;
   wire n_5_4494;
   wire n_5_4540;
   wire n_5_4541;
   wire n_5_4544;
   wire n_5_4545;
   wire n_5_4546;
   wire n_5_4547;
   wire n_5_4550;
   wire n_5_4556;
   wire n_5_4599;
   wire n_5_4603;
   wire n_5_3891;
   wire n_5_3946;
   wire n_5_4769;
   wire n_5_3947;
   wire n_5_4772;
   wire n_5_4773;
   wire n_5_4796;
   wire n_5_650;
   wire n_5_240;
   wire n_5_4797;
   wire n_5_4798;
   wire n_5_4799;
   wire n_5_4800;
   wire n_5_4542;
   wire n_5_4801;
   wire n_5_3955;
   wire n_5_4803;
   wire n_5_3966;
   wire n_5_3974;
   wire n_5_3978;
   wire n_5_3995;
   wire n_5_4307;
   wire n_5_4310;
   wire n_5_4344;
   wire n_5_4345;
   wire n_5_4349;
   wire n_5_4372;
   wire n_5_4459;
   wire n_5_4491;
   wire n_5_4502;
   wire n_5_4521;
   wire n_5_4523;
   wire n_5_4555;
   wire n_5_4567;
   wire n_5_4571;
   wire n_5_4572;
   wire n_5_4594;
   wire n_5_4604;
   wire n_5_4605;
   wire n_5_4608;
   wire n_5_4615;
   wire n_5_4616;
   wire n_5_4624;
   wire n_5_4641;
   wire n_5_4669;
   wire n_5_4710;
   wire n_5_4720;
   wire n_5_4721;
   wire n_5_4724;
   wire n_5_4726;
   wire n_5_4727;
   wire n_5_4733;
   wire n_5_4735;
   wire n_5_4770;
   wire n_5_4771;
   wire n_5_4802;
   wire n_5_4804;
   wire n_5_4805;
   wire n_5_4806;
   wire n_5_204;
   wire n_5_3862;
   wire n_5_4807;
   wire n_5_4808;
   wire n_5_4809;
   wire n_5_4810;
   wire n_5_4811;
   wire n_5_4812;
   wire n_5_4813;
   wire n_5_4814;
   wire n_7_0;
   wire n_7_1;
   wire n_7_2;
   wire n_7_3;
   wire n_7_4;
   wire n_7_5;
   wire n_7_6;
   wire n_7_7;
   wire n_7_8;
   wire n_7_9;
   wire n_7_10;
   wire n_7_11;
   wire n_7_12;
   wire n_7_13;
   wire n_7_14;
   wire n_7_15;
   wire n_7_16;
   wire n_7_17;
   wire n_7_19;
   wire n_7_21;
   wire n_7_22;
   wire n_7_20;
   wire n_7_24;
   wire n_7_23;
   wire n_7_26;
   wire n_7_27;
   wire n_7_28;
   wire n_7_29;
   wire n_7_30;
   wire n_7_31;
   wire n_7_32;
   wire n_7_33;
   wire n_7_34;
   wire n_7_35;
   wire n_7_36;
   wire n_7_37;
   wire n_7_38;
   wire n_7_39;
   wire n_7_40;
   wire n_7_41;
   wire n_7_42;
   wire n_7_43;
   wire n_7_44;
   wire n_7_45;
   wire n_7_46;
   wire n_7_47;
   wire n_7_48;
   wire n_7_49;
   wire n_7_50;
   wire n_7_51;
   wire n_7_52;
   wire n_7_53;
   wire n_7_54;
   wire n_7_55;
   wire n_7_56;
   wire n_7_57;
   wire n_7_58;
   wire n_7_59;
   wire n_7_60;
   wire n_7_61;
   wire n_7_62;
   wire n_7_63;
   wire n_7_64;
   wire n_7_65;
   wire n_7_66;
   wire n_7_67;
   wire n_7_68;
   wire n_7_69;
   wire n_7_70;
   wire n_7_71;
   wire n_7_72;
   wire n_7_73;
   wire n_7_74;
   wire n_7_75;
   wire n_7_76;
   wire n_7_77;
   wire n_7_78;
   wire n_7_79;
   wire n_7_80;
   wire n_7_81;
   wire n_7_82;
   wire n_7_83;
   wire n_7_84;
   wire n_7_85;
   wire n_7_86;
   wire n_7_87;
   wire n_7_88;
   wire n_7_89;
   wire n_7_90;
   wire n_7_91;
   wire n_7_92;
   wire n_7_93;
   wire n_7_94;
   wire n_7_95;
   wire n_7_96;
   wire n_7_97;
   wire n_7_98;
   wire n_7_99;
   wire n_7_100;
   wire n_7_101;
   wire n_7_102;
   wire n_7_103;
   wire n_7_104;
   wire n_7_105;
   wire n_7_106;
   wire n_7_107;
   wire n_7_108;
   wire n_7_109;
   wire n_7_110;
   wire n_7_111;
   wire n_7_112;
   wire n_7_113;
   wire n_7_114;
   wire n_7_115;
   wire n_7_116;
   wire n_7_117;
   wire n_7_118;
   wire n_7_119;
   wire n_7_120;
   wire n_7_176;
   wire n_7_18;
   wire n_7_177;
   wire n_7_25;
   wire n_7_121;
   wire n_7_178;
   wire n_7_122;
   wire n_7_179;
   wire n_7_123;
   wire n_7_180;
   wire n_7_181;
   wire n_7_124;
   wire n_7_182;
   wire n_7_125;
   wire n_7_126;
   wire n_7_127;
   wire n_7_128;
   wire n_7_129;
   wire n_7_130;
   wire n_7_131;
   wire n_7_133;
   wire n_7_138;
   wire n_7_132;
   wire n_7_142;
   wire n_7_183;
   wire n_7_184;
   wire n_7_144;
   wire n_7_145;
   wire n_7_146;
   wire n_7_147;
   wire n_7_185;
   wire n_7_135;
   wire n_7_150;
   wire n_7_151;
   wire n_7_152;
   wire n_7_186;
   wire n_7_153;
   wire n_7_154;
   wire n_7_155;
   wire n_7_156;
   wire n_7_157;
   wire n_7_158;
   wire n_7_159;
   wire n_7_160;
   wire n_7_161;
   wire n_7_162;
   wire n_7_164;
   wire n_7_165;
   wire n_7_166;
   wire n_7_167;
   wire n_7_168;
   wire n_7_169;
   wire n_7_187;
   wire n_7_170;
   wire n_7_171;
   wire n_7_172;
   wire n_7_173;
   wire n_7_174;
   wire n_7_188;
   wire n_7_189;
   wire n_7_190;
   wire n_7_191;
   wire n_7_136;
   wire n_7_194;
   wire n_7_195;
   wire n_7_137;
   wire n_7_139;
   wire n_7_140;
   wire n_7_143;
   wire n_7_148;
   wire n_7_149;
   wire n_7_134;
   wire n_7_175;
   wire n_7_192;
   wire n_7_193;
   wire n_7_141;
   wire n_7_197;
   wire n_7_198;
   wire n_7_200;
   wire n_7_204;
   wire n_7_205;
   wire n_7_201;
   wire n_7_202;
   wire n_7_203;
   wire n_7_163;
   wire n_7_196;
   wire n_7_199;
   wire n_7_206;
   wire n_7_207;
   wire n_7_208;
   wire n_8_0;
   wire n_8_1;
   wire n_8_410;
   wire n_8_3;
   wire n_8_7;
   wire n_8_20;
   wire n_8_21;
   wire n_8_23;
   wire n_8_26;
   wire n_8_36;
   wire n_8_8;
   wire n_8_12;
   wire n_8_411;
   wire n_8_412;
   wire n_8_413;
   wire n_8_414;
   wire n_8_65;
   wire n_8_67;
   wire n_8_35;
   wire n_8_49;
   wire n_8_54;
   wire n_8_31;
   wire n_8_70;
   wire n_8_71;
   wire n_8_72;
   wire n_8_76;
   wire n_8_77;
   wire n_8_79;
   wire n_8_80;
   wire n_8_415;
   wire n_8_27;
   wire n_8_28;
   wire n_8_56;
   wire n_8_24;
   wire n_8_82;
   wire n_8_83;
   wire n_8_416;
   wire n_8_2;
   wire n_8_25;
   wire n_8_32;
   wire n_8_44;
   wire n_8_46;
   wire n_8_47;
   wire n_8_48;
   wire n_8_57;
   wire n_8_417;
   wire n_8_418;
   wire n_8_419;
   wire n_8_88;
   wire n_8_43;
   wire n_8_45;
   wire n_8_53;
   wire n_8_58;
   wire n_8_81;
   wire n_8_60;
   wire n_8_61;
   wire n_8_64;
   wire n_8_66;
   wire n_8_73;
   wire n_8_75;
   wire n_8_86;
   wire n_8_87;
   wire n_8_420;
   wire n_8_421;
   wire n_8_9;
   wire n_8_13;
   wire n_8_38;
   wire n_8_39;
   wire n_8_4;
   wire n_8_5;
   wire n_8_17;
   wire n_8_18;
   wire n_8_11;
   wire n_8_40;
   wire n_8_19;
   wire n_8_6;
   wire n_8_10;
   wire n_8_14;
   wire n_8_15;
   wire n_8_16;
   wire n_8_22;
   wire n_8_29;
   wire n_8_30;
   wire n_8_33;
   wire n_8_34;
   wire n_8_37;
   wire n_8_41;
   wire n_8_42;
   wire n_8_422;
   wire n_8_63;
   wire n_8_50;
   wire n_8_51;
   wire n_8_52;
   wire n_8_182;
   wire n_8_55;
   wire n_8_59;
   wire n_8_62;
   wire n_8_68;
   wire n_8_69;
   wire n_8_74;
   wire n_8_78;
   wire n_8_84;
   wire n_8_85;
   wire n_8_89;
   wire n_8_90;
   wire n_8_91;
   wire n_8_92;
   wire n_8_93;
   wire n_8_94;
   wire n_8_95;
   wire n_8_96;
   wire n_8_97;
   wire n_8_98;
   wire n_8_99;
   wire n_8_100;
   wire n_8_101;
   wire n_8_102;
   wire n_8_103;
   wire n_8_104;
   wire n_8_105;
   wire n_8_106;
   wire n_8_107;
   wire n_8_108;
   wire n_8_183;
   wire n_8_109;
   wire n_8_110;
   wire n_8_111;
   wire n_8_112;
   wire n_8_113;
   wire n_8_114;
   wire n_8_115;
   wire n_8_116;
   wire n_8_117;
   wire n_8_118;
   wire n_8_119;
   wire n_8_120;
   wire n_8_423;
   wire n_8_290;
   wire n_8_292;
   wire n_8_121;
   wire n_8_122;
   wire n_8_424;
   wire n_8_425;
   wire n_8_123;
   wire n_8_124;
   wire n_8_426;
   wire n_8_427;
   wire n_8_428;
   wire n_8_429;
   wire n_8_430;
   wire n_8_431;
   wire n_8_432;
   wire n_8_125;
   wire n_8_126;
   wire n_8_433;
   wire n_8_434;
   wire n_8_127;
   wire n_8_435;
   wire n_8_436;
   wire n_8_437;
   wire n_8_128;
   wire n_8_129;
   wire n_8_130;
   wire n_8_131;
   wire n_8_132;
   wire n_8_133;
   wire n_8_134;
   wire n_8_135;
   wire n_8_438;
   wire n_8_136;
   wire n_8_137;
   wire n_8_138;
   wire n_8_439;
   wire n_8_139;
   wire n_8_140;
   wire n_8_141;
   wire n_8_142;
   wire n_8_143;
   wire n_8_144;
   wire n_8_145;
   wire n_8_192;
   wire n_8_146;
   wire n_8_147;
   wire n_8_148;
   wire n_8_149;
   wire n_8_150;
   wire n_8_151;
   wire n_8_152;
   wire n_8_153;
   wire n_8_154;
   wire n_8_155;
   wire n_8_156;
   wire n_8_157;
   wire n_8_158;
   wire n_8_159;
   wire n_8_160;
   wire n_8_161;
   wire n_8_162;
   wire n_8_163;
   wire n_8_164;
   wire n_8_165;
   wire n_8_166;
   wire n_8_167;
   wire n_8_168;
   wire n_8_169;
   wire n_8_170;
   wire n_8_171;
   wire n_8_172;
   wire n_8_173;
   wire n_8_174;
   wire n_8_175;
   wire n_8_193;
   wire n_8_176;
   wire n_8_177;
   wire n_8_440;
   wire n_8_441;
   wire n_8_178;
   wire n_8_179;
   wire n_8_180;
   wire n_8_181;
   wire n_8_184;
   wire n_8_185;
   wire n_8_186;
   wire n_8_187;
   wire n_8_442;
   wire n_8_188;
   wire n_8_189;
   wire n_8_190;
   wire n_8_191;
   wire n_8_194;
   wire n_8_195;
   wire n_8_196;
   wire n_8_443;
   wire n_8_197;
   wire n_8_444;
   wire n_8_198;
   wire n_8_199;
   wire n_8_200;
   wire n_8_201;
   wire n_8_445;
   wire n_8_202;
   wire n_8_203;
   wire n_8_204;
   wire n_8_205;
   wire n_8_206;
   wire n_8_207;
   wire n_8_208;
   wire n_8_209;
   wire n_8_210;
   wire n_8_211;
   wire n_8_212;
   wire n_8_294;
   wire n_8_213;
   wire n_8_214;
   wire n_8_215;
   wire n_8_295;
   wire n_8_216;
   wire n_8_217;
   wire n_8_218;
   wire n_8_219;
   wire n_8_220;
   wire n_8_221;
   wire n_8_222;
   wire n_8_223;
   wire n_8_224;
   wire n_8_225;
   wire n_8_298;
   wire n_8_226;
   wire n_8_227;
   wire n_8_228;
   wire n_8_229;
   wire n_8_230;
   wire n_8_231;
   wire n_8_232;
   wire n_8_233;
   wire n_8_234;
   wire n_8_235;
   wire n_8_236;
   wire n_8_237;
   wire n_8_238;
   wire n_8_239;
   wire n_8_240;
   wire n_8_241;
   wire n_8_242;
   wire n_8_243;
   wire n_8_244;
   wire n_8_245;
   wire n_8_246;
   wire n_8_446;
   wire n_8_447;
   wire n_8_247;
   wire n_8_248;
   wire n_8_249;
   wire n_8_250;
   wire n_8_251;
   wire n_8_448;
   wire n_8_300;
   wire n_8_254;
   wire n_8_255;
   wire n_8_449;
   wire n_8_450;
   wire n_8_258;
   wire n_8_259;
   wire n_8_260;
   wire n_8_261;
   wire n_8_263;
   wire n_8_264;
   wire n_8_451;
   wire n_8_266;
   wire n_8_267;
   wire n_8_268;
   wire n_8_269;
   wire n_8_271;
   wire n_8_272;
   wire n_8_273;
   wire n_8_302;
   wire n_8_274;
   wire n_8_275;
   wire n_8_276;
   wire n_8_452;
   wire n_8_304;
   wire n_8_277;
   wire n_8_453;
   wire n_8_281;
   wire n_8_454;
   wire n_8_283;
   wire n_8_284;
   wire n_8_455;
   wire n_8_286;
   wire n_8_287;
   wire n_8_288;
   wire n_8_289;
   wire n_8_456;
   wire n_8_308;
   wire n_8_309;
   wire n_8_310;
   wire n_8_311;
   wire n_8_312;
   wire n_8_252;
   wire n_8_253;
   wire n_8_313;
   wire n_8_457;
   wire n_8_458;
   wire n_8_459;
   wire n_8_460;
   wire n_8_461;
   wire n_8_462;
   wire n_8_463;
   wire n_8_464;
   wire n_8_465;
   wire n_8_466;
   wire n_8_467;
   wire n_8_468;
   wire n_8_469;
   wire n_8_470;
   wire n_8_471;
   wire n_8_472;
   wire n_8_473;
   wire n_8_474;
   wire n_8_475;
   wire n_8_476;
   wire n_8_477;
   wire n_8_478;
   wire n_8_479;
   wire n_8_480;
   wire n_8_481;
   wire n_8_482;
   wire n_8_483;
   wire n_8_256;
   wire n_8_257;
   wire n_8_262;
   wire n_8_265;
   wire n_8_270;
   wire n_8_278;
   wire n_8_279;
   wire n_8_280;
   wire n_8_484;
   wire n_8_282;
   wire n_8_285;
   wire n_8_291;
   wire n_8_485;
   wire n_8_293;
   wire n_8_296;
   wire n_8_486;
   wire n_8_487;
   wire n_8_488;
   wire n_8_489;
   wire n_8_490;
   wire n_8_491;
   wire n_8_492;
   wire n_8_297;
   wire n_8_299;
   wire n_8_301;
   wire n_8_493;
   wire n_8_303;
   wire n_8_305;
   wire n_8_306;
   wire n_8_307;
   wire n_8_494;
   wire n_8_495;
   wire n_8_496;
   wire n_8_497;
   wire n_8_498;
   wire n_8_499;
   wire n_8_500;
   wire n_8_501;
   wire n_8_502;
   wire n_8_503;
   wire n_8_314;
   wire n_8_315;
   wire n_8_316;
   wire n_8_317;
   wire n_8_318;
   wire n_8_319;
   wire n_8_320;
   wire n_8_321;
   wire n_8_504;
   wire n_8_322;
   wire n_8_323;
   wire n_8_324;
   wire n_8_325;
   wire n_8_326;
   wire n_8_327;
   wire n_8_328;
   wire n_8_329;
   wire n_8_330;
   wire n_8_331;
   wire n_8_332;
   wire n_8_333;
   wire n_8_505;
   wire n_8_334;
   wire n_8_335;
   wire n_8_336;
   wire n_8_337;
   wire n_8_338;
   wire n_8_339;
   wire n_8_340;
   wire n_8_341;
   wire n_8_342;
   wire n_8_343;
   wire n_8_344;
   wire n_8_345;
   wire n_8_346;
   wire n_8_347;
   wire n_8_348;
   wire n_8_349;
   wire n_8_350;
   wire n_8_351;
   wire n_8_352;
   wire n_8_353;
   wire n_8_354;
   wire n_8_355;
   wire n_8_356;
   wire n_8_357;
   wire n_8_358;
   wire n_8_359;
   wire n_8_360;
   wire n_8_361;
   wire n_8_362;
   wire n_8_363;
   wire n_8_364;
   wire n_8_365;
   wire n_8_366;
   wire n_8_367;
   wire n_8_368;
   wire n_8_369;
   wire n_8_370;
   wire n_8_371;
   wire n_8_372;
   wire n_8_373;
   wire n_8_374;
   wire n_8_375;
   wire n_8_376;
   wire n_8_377;
   wire n_8_378;
   wire n_8_379;
   wire n_8_380;
   wire n_8_381;
   wire n_8_382;
   wire n_8_383;
   wire n_8_384;
   wire n_8_385;
   wire n_8_506;
   wire n_8_386;
   wire n_8_387;
   wire n_8_388;
   wire n_8_389;
   wire n_8_390;
   wire n_8_391;
   wire n_8_392;
   wire n_8_507;
   wire n_8_393;
   wire n_8_394;
   wire n_8_395;
   wire n_8_396;
   wire n_8_397;
   wire n_8_398;
   wire n_8_399;
   wire n_8_400;
   wire n_8_401;
   wire n_8_402;
   wire n_8_403;
   wire n_8_508;
   wire n_8_404;
   wire n_8_405;
   wire n_8_406;
   wire n_8_407;
   wire n_8_408;
   wire n_8_409;
   wire n_8_509;
   wire n_8_510;
   wire n_8_511;
   wire n_8_512;
   wire n_8_513;
   wire n_8_514;
   wire n_8_515;
   wire n_8_516;
   wire n_8_517;
   wire n_8_518;
   wire n_8_519;
   wire n_8_520;
   wire n_8_521;
   wire n_8_522;
   wire n_8_523;
   wire n_8_524;
   wire n_8_525;
   wire n_8_526;
   wire n_8_527;
   wire n_8_528;
   wire n_8_529;
   wire n_8_530;
   wire n_8_531;
   wire n_8_532;
   wire n_8_533;
   wire n_8_534;
   wire n_8_535;
   wire n_8_536;
   wire n_8_537;
   wire n_8_538;
   wire n_8_539;
   wire n_8_540;
   wire n_8_541;
   wire n_8_542;
   wire n_8_543;
   wire n_8_544;
   wire n_8_545;
   wire n_8_546;
   wire n_8_547;
   wire n_8_548;
   wire n_8_549;
   wire n_8_550;
   wire n_8_551;
   wire n_8_552;
   wire n_8_553;
   wire n_8_554;
   wire n_8_555;
   wire n_8_556;
   wire n_8_557;
   wire n_8_558;
   wire n_8_559;
   wire n_8_560;
   wire n_8_561;
   wire n_8_562;
   wire n_8_563;
   wire n_8_564;
   wire n_8_565;
   wire n_8_566;
   wire n_8_567;
   wire n_8_568;
   wire n_8_569;
   wire n_8_570;
   wire n_8_571;
   wire n_8_572;
   wire n_8_573;
   wire n_8_574;
   wire n_8_575;
   wire n_8_576;
   wire n_8_577;
   wire n_8_578;
   wire n_8_579;
   wire n_8_580;
   wire n_8_581;
   wire n_8_582;
   wire n_8_583;
   wire n_8_584;
   wire n_8_585;
   wire n_8_586;
   wire n_8_587;
   wire n_8_588;
   wire n_8_589;
   wire n_8_590;
   wire n_8_591;
   wire n_8_592;

   datapath__2_486 i_1 (.R({uc_0, uc_1, uc_2, uc_3, n_76, n_73, n_55, n_60, n_69, 
      n_68, n_66, n_58, n_65, n_59, n_56, m[0], uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, 
      uc_20}), .L({uc_21, uc_22, uc_23, uc_24, n_86, n_92, n_85, n_84, n_91, 
      n_90, n_83, n_82, n_81, n_93, n_80, n_79, uc_25, uc_26, uc_27, uc_28, 
      uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, 
      uc_39, uc_40, uc_41}), .plus({uc_42, uc_43, uc_44, uc_45, n_11, n_10, n_9, 
      n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_46, uc_47, uc_48, uc_49, 
      uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, 
      uc_60, uc_61, uc_62}));
   NAND2_X1 i_2_0 (.A1(n_102), .A2(n_2_32), .ZN(n_2_0));
   NAND2_X1 i_2_1 (.A1(n_112), .A2(n_2_30), .ZN(n_2_1));
   NAND2_X1 i_2_2 (.A1(n_125), .A2(n_2_34), .ZN(n_2_2));
   NAND3_X1 i_2_3 (.A1(n_2_0), .A2(n_2_1), .A3(n_2_2), .ZN(n_12));
   NAND2_X1 i_2_4 (.A1(n_113), .A2(n_2_30), .ZN(n_2_3));
   NAND2_X1 i_2_5 (.A1(n_103), .A2(n_2_32), .ZN(n_2_4));
   NAND2_X1 i_2_6 (.A1(n_123), .A2(n_2_34), .ZN(n_2_5));
   NAND3_X1 i_2_7 (.A1(n_2_3), .A2(n_2_4), .A3(n_2_5), .ZN(n_13));
   NAND2_X1 i_2_8 (.A1(n_108), .A2(n_2_32), .ZN(n_2_6));
   NAND2_X1 i_2_9 (.A1(n_122), .A2(n_2_34), .ZN(n_2_7));
   INV_X1 i_2_10 (.A(n_2_7), .ZN(n_2_8));
   AOI21_X1 i_2_11 (.A(n_2_8), .B1(n_117), .B2(n_2_30), .ZN(n_2_9));
   NAND2_X1 i_2_12 (.A1(n_2_6), .A2(n_2_9), .ZN(n_14));
   NAND2_X1 i_2_13 (.A1(n_116), .A2(n_2_30), .ZN(n_2_10));
   NAND2_X1 i_2_14 (.A1(n_105), .A2(n_2_32), .ZN(n_2_11));
   NAND2_X1 i_2_15 (.A1(n_128), .A2(n_2_34), .ZN(n_2_12));
   NAND3_X1 i_2_16 (.A1(n_2_10), .A2(n_2_11), .A3(n_2_12), .ZN(n_15));
   NAND2_X1 i_2_17 (.A1(n_120), .A2(n_2_30), .ZN(n_2_13));
   NAND2_X1 i_2_18 (.A1(n_110), .A2(n_2_32), .ZN(n_2_14));
   NAND2_X1 i_2_19 (.A1(n_130), .A2(n_2_34), .ZN(n_2_15));
   NAND3_X1 i_2_20 (.A1(n_2_13), .A2(n_2_14), .A3(n_2_15), .ZN(n_16));
   NAND2_X1 i_2_21 (.A1(n_109), .A2(n_2_32), .ZN(n_2_16));
   NAND2_X1 i_2_22 (.A1(n_118), .A2(n_2_30), .ZN(n_2_17));
   NAND2_X1 i_2_23 (.A1(n_131), .A2(n_2_34), .ZN(n_2_18));
   NAND3_X1 i_2_24 (.A1(n_2_16), .A2(n_2_17), .A3(n_2_18), .ZN(n_17));
   NAND2_X1 i_2_25 (.A1(n_124), .A2(n_2_30), .ZN(n_2_19));
   NAND2_X1 i_2_26 (.A1(n_111), .A2(n_2_32), .ZN(n_2_20));
   NAND2_X1 i_2_27 (.A1(n_133), .A2(n_2_34), .ZN(n_2_21));
   NAND3_X1 i_2_28 (.A1(n_2_19), .A2(n_2_20), .A3(n_2_21), .ZN(n_18));
   NAND2_X1 i_2_29 (.A1(n_114), .A2(n_2_30), .ZN(n_2_22));
   NAND2_X1 i_2_30 (.A1(n_106), .A2(n_2_32), .ZN(n_2_23));
   NAND2_X1 i_2_31 (.A1(n_129), .A2(n_2_34), .ZN(n_2_24));
   NAND3_X1 i_2_32 (.A1(n_2_22), .A2(n_2_23), .A3(n_2_24), .ZN(n_19));
   NAND2_X1 i_2_33 (.A1(n_104), .A2(n_2_32), .ZN(n_2_25));
   NAND2_X1 i_2_34 (.A1(n_115), .A2(n_2_30), .ZN(n_2_26));
   NAND2_X1 i_2_35 (.A1(n_132), .A2(n_2_34), .ZN(n_2_27));
   NAND3_X1 i_2_36 (.A1(n_2_25), .A2(n_2_26), .A3(n_2_27), .ZN(n_20));
   INV_X1 i_2_37 (.A(r[12]), .ZN(n_2_28));
   NAND2_X1 i_2_38 (.A1(r[13]), .A2(n_2_28), .ZN(n_2_29));
   INV_X1 i_2_39 (.A(n_2_29), .ZN(n_2_30));
   NAND2_X1 i_2_40 (.A1(n_119), .A2(n_2_30), .ZN(n_2_31));
   NOR2_X1 i_2_41 (.A1(r[13]), .A2(n_2_28), .ZN(n_2_32));
   NAND2_X1 i_2_42 (.A1(n_107), .A2(n_2_32), .ZN(n_2_33));
   XNOR2_X1 i_2_43 (.A(r[13]), .B(r[12]), .ZN(n_2_34));
   NAND2_X1 i_2_44 (.A1(n_126), .A2(n_2_34), .ZN(n_2_35));
   NAND3_X1 i_2_45 (.A1(n_2_31), .A2(n_2_33), .A3(n_2_35), .ZN(n_21));
   datapath__2_495 i_4 (.R({uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, 
      n_60, n_69, n_68, n_66, n_58, n_65, n_59, n_56, m[0], uc_70, uc_71, uc_72, 
      uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, 
      uc_83, uc_84, uc_85, uc_86}), .L({uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, 
      uc_93, n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, uc_94, uc_95, 
      uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, 
      uc_106, uc_107, uc_108, uc_109, uc_110}), .plus({uc_111, uc_112, uc_113, 
      uc_114, uc_115, uc_116, uc_117, n_30, n_29, n_28, n_27, n_26, n_25, n_24, 
      n_23, n_22, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, uc_124, uc_125, 
      uc_126, uc_127, uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, uc_134}));
   datapath__2_498 i_6 (.R({uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, 
      uc_141, uc_142, n_69, n_68, n_66, n_58, n_65, n_59, n_56, m[0], uc_143, 
      uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, 
      uc_153, uc_154, uc_155, uc_156, uc_157, uc_158, uc_159}), .L({uc_160, 
      uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, n_100, n_101, n_99, 
      n_98, n_97, n_96, n_95, n_94, uc_168, uc_169, uc_170, uc_171, uc_172, 
      uc_173, uc_174, uc_175, uc_176, uc_177, uc_178, uc_179, uc_180, uc_181, 
      uc_182, uc_183, uc_184}), .plus({uc_185, uc_186, uc_187, uc_188, uc_189, 
      uc_190, uc_191, uc_192, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, 
      uc_193, uc_194, uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, 
      uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, uc_208, uc_209}));
   datapath__2_752 i_3 (.R({uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, 
      uc_216, uc_217, m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_218, 
      uc_219, uc_220, uc_221, uc_222, uc_223, uc_224, uc_225, uc_226, uc_227, 
      uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, uc_234}), .L({uc_235, 
      uc_236, uc_237, uc_238, uc_239, uc_240, uc_241, uc_242, n_100, n_101, n_99, 
      n_98, n_97, n_96, n_95, n_94, uc_243, uc_244, uc_245, uc_246, uc_247, 
      uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, uc_254, uc_255, uc_256, 
      uc_257, uc_258, uc_259}), .plus({uc_260, uc_261, uc_262, uc_263, uc_264, 
      uc_265, uc_266, uc_267, n_46, n_45, n_44, n_43, n_42, n_41, n_40, n_39, 
      uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, 
      uc_277, uc_278, uc_279, uc_280, uc_281, uc_282, uc_283, uc_284}));
   NOR4_X1 i_45_0 (.A1(r[0]), .A2(r[1]), .A3(r[2]), .A4(r[3]), .ZN(n_45_0));
   NOR4_X1 i_45_1 (.A1(r[4]), .A2(r[5]), .A3(r[6]), .A4(r[7]), .ZN(n_45_1));
   NOR4_X1 i_45_2 (.A1(r[8]), .A2(r[9]), .A3(r[10]), .A4(r[11]), .ZN(n_45_2));
   NOR4_X1 i_45_3 (.A1(r[12]), .A2(r[13]), .A3(r[14]), .A4(r[15]), .ZN(n_45_3));
   NAND4_X1 i_45_4 (.A1(n_45_0), .A2(n_45_1), .A3(n_45_2), .A4(n_45_3), .ZN(
      n_45_4));
   NOR4_X1 i_45_5 (.A1(m[0]), .A2(m[1]), .A3(m[2]), .A4(m[3]), .ZN(n_45_5));
   NOR4_X1 i_45_6 (.A1(m[4]), .A2(m[5]), .A3(m[6]), .A4(m[7]), .ZN(n_45_6));
   NOR4_X1 i_45_7 (.A1(m[8]), .A2(m[9]), .A3(m[10]), .A4(m[11]), .ZN(n_45_7));
   NOR4_X1 i_45_8 (.A1(m[12]), .A2(m[13]), .A3(m[14]), .A4(m[15]), .ZN(n_45_8));
   NAND4_X1 i_45_9 (.A1(n_45_5), .A2(n_45_6), .A3(n_45_7), .A4(n_45_8), .ZN(
      n_45_9));
   AND2_X1 i_45_10 (.A1(n_45_9), .A2(n_45_4), .ZN(n_47));
   NAND2_X1 i_0_16 (.A1(n_55), .A2(n_0_3), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_48));
   NAND2_X1 i_0_4 (.A1(n_75), .A2(n_0_3), .ZN(n_0_11));
   INV_X1 i_0_6 (.A(n_0_11), .ZN(n_49));
   NAND2_X1 i_0_7 (.A1(n_0_89), .A2(n_0_3), .ZN(n_0_12));
   INV_X1 i_0_13 (.A(n_0_12), .ZN(n_50));
   NAND2_X1 i_0_26 (.A1(n_53), .A2(n_0_3), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(n_51));
   NAND2_X1 i_0_28 (.A1(n_54), .A2(n_0_3), .ZN(n_0_14));
   INV_X1 i_0_29 (.A(n_0_14), .ZN(n_52));
   AOI21_X1 i_0_36 (.A(n_0_5), .B1(m[14]), .B2(n_0_196), .ZN(n_53));
   XNOR2_X1 i_0_39 (.A(m[15]), .B(n_0_5), .ZN(n_54));
   NOR4_X1 i_0_40 (.A1(m[13]), .A2(m[12]), .A3(m[14]), .A4(n_0_9), .ZN(n_0_5));
   INV_X1 i_0_45 (.A(n_0_1), .ZN(n_55));
   NAND2_X1 i_0_46 (.A1(n_0_2), .A2(n_0_159), .ZN(n_0_1));
   NAND2_X1 i_0_47 (.A1(n_0_111), .A2(m[9]), .ZN(n_0_2));
   OAI21_X1 i_0_12 (.A(n_0_71), .B1(n_0_122), .B2(n_0_18), .ZN(n_0_7));
   INV_X1 i_0_52 (.A(m[9]), .ZN(n_0_20));
   INV_X1 i_0_55 (.A(m[10]), .ZN(n_0_18));
   XNOR2_X1 i_0_5 (.A(m[1]), .B(m[0]), .ZN(n_0_21));
   INV_X1 i_0_107 (.A(m[8]), .ZN(n_0_24));
   INV_X1 i_0_2 (.A(m[0]), .ZN(n_0_28));
   INV_X1 i_0_8 (.A(n_0_21), .ZN(n_56));
   INV_X1 i_0_0 (.A(r[0]), .ZN(n_0_29));
   NOR2_X1 i_0_9 (.A1(n_0_21), .A2(n_0_29), .ZN(n_57));
   NAND4_X1 i_0_20 (.A1(n_0_31), .A2(n_0_32), .A3(n_0_33), .A4(n_0_34), .ZN(
      n_0_0));
   INV_X1 i_0_53 (.A(m[6]), .ZN(n_0_31));
   INV_X1 i_0_86 (.A(m[7]), .ZN(n_0_32));
   INV_X1 i_0_87 (.A(m[5]), .ZN(n_0_33));
   INV_X1 i_0_89 (.A(m[4]), .ZN(n_0_34));
   NOR2_X1 i_0_129 (.A1(m[6]), .A2(m[7]), .ZN(n_0_36));
   NOR2_X1 i_0_130 (.A1(m[5]), .A2(m[0]), .ZN(n_0_37));
   NOR2_X1 i_0_131 (.A1(m[4]), .A2(m[1]), .ZN(n_0_38));
   NOR2_X1 i_0_132 (.A1(m[2]), .A2(m[3]), .ZN(n_0_39));
   NAND4_X1 i_0_133 (.A1(n_0_36), .A2(n_0_37), .A3(n_0_38), .A4(n_0_39), 
      .ZN(n_0_40));
   INV_X1 i_0_104 (.A(n_0_108), .ZN(n_58));
   INV_X1 i_0_14 (.A(n_0_35), .ZN(n_59));
   NAND2_X1 i_0_1 (.A1(n_0_132), .A2(n_0_133), .ZN(n_0_35));
   INV_X1 i_0_11 (.A(m[7]), .ZN(n_0_42));
   INV_X1 i_0_76 (.A(m[7]), .ZN(n_0_43));
   NAND3_X1 i_0_60 (.A1(n_0_43), .A2(n_0_186), .A3(n_0_185), .ZN(n_0_46));
   INV_X1 i_0_70 (.A(n_0_46), .ZN(n_0_47));
   INV_X1 i_0_128 (.A(m[6]), .ZN(n_0_49));
   INV_X1 i_0_134 (.A(m[5]), .ZN(n_0_50));
   INV_X1 i_0_148 (.A(m[0]), .ZN(n_0_51));
   NAND3_X1 i_0_110 (.A1(n_0_49), .A2(n_0_50), .A3(n_0_51), .ZN(n_0_52));
   INV_X1 i_0_72 (.A(n_0_52), .ZN(n_0_53));
   BUF_X1 rt_shieldBuf__2__2__0 (.A(r[0]), .Z(n_0_3));
   INV_X1 i_0_137 (.A(m[4]), .ZN(n_0_55));
   INV_X1 i_0_149 (.A(m[3]), .ZN(n_0_56));
   INV_X1 i_0_150 (.A(m[8]), .ZN(n_0_57));
   NAND3_X1 i_0_151 (.A1(n_0_55), .A2(n_0_56), .A3(n_0_57), .ZN(n_0_58));
   INV_X1 i_0_74 (.A(n_0_58), .ZN(n_0_59));
   INV_X1 i_0_116 (.A(n_0_114), .ZN(n_60));
   INV_X1 i_0_22 (.A(r[0]), .ZN(n_0_60));
   INV_X1 i_0_19 (.A(m[6]), .ZN(n_0_26));
   INV_X1 i_0_25 (.A(m[5]), .ZN(n_0_15));
   INV_X1 i_0_34 (.A(m[0]), .ZN(n_0_22));
   INV_X1 i_0_44 (.A(m[4]), .ZN(n_0_41));
   INV_X1 i_0_146 (.A(m[0]), .ZN(n_0_65));
   INV_X1 i_0_147 (.A(m[2]), .ZN(n_0_66));
   INV_X1 i_0_157 (.A(m[1]), .ZN(n_0_67));
   INV_X1 i_0_158 (.A(m[3]), .ZN(n_0_68));
   INV_X1 i_0_156 (.A(n_0_100), .ZN(n_0_74));
   NAND2_X1 i_0_162 (.A1(n_0_80), .A2(n_0_74), .ZN(n_0_75));
   NOR2_X1 i_0_142 (.A1(m[12]), .A2(n_0_9), .ZN(n_0_77));
   INV_X1 i_0_160 (.A(n_0_201), .ZN(n_0_9));
   INV_X1 i_0_167 (.A(m[13]), .ZN(n_0_84));
   INV_X1 i_0_168 (.A(m[12]), .ZN(n_0_85));
   NAND2_X1 i_0_169 (.A1(n_0_84), .A2(n_0_85), .ZN(n_0_86));
   NOR2_X1 i_0_170 (.A1(n_0_9), .A2(n_0_86), .ZN(n_0_87));
   INV_X1 i_0_171 (.A(n_0_77), .ZN(n_0_88));
   AOI21_X1 i_0_172 (.A(n_0_87), .B1(n_0_88), .B2(m[13]), .ZN(n_0_89));
   INV_X1 i_0_117 (.A(m[0]), .ZN(n_0_23));
   INV_X1 i_0_139 (.A(m[5]), .ZN(n_0_27));
   NAND4_X1 i_0_18 (.A1(n_0_42), .A2(n_0_63), .A3(n_0_64), .A4(n_0_72), .ZN(
      n_0_93));
   NAND2_X1 i_0_49 (.A1(n_0_26), .A2(n_0_42), .ZN(n_0_97));
   INV_X1 i_0_50 (.A(n_0_97), .ZN(n_0_98));
   BUF_X1 rt_shieldBuf__2__2__1 (.A(n_0_89), .Z(n_61));
   INV_X1 i_0_79 (.A(m[4]), .ZN(n_0_44));
   INV_X1 i_0_95 (.A(m[1]), .ZN(n_0_61));
   INV_X1 i_0_96 (.A(m[3]), .ZN(n_0_62));
   NAND2_X1 i_0_73 (.A1(n_0_130), .A2(n_0_105), .ZN(n_0_108));
   NAND3_X1 i_0_114 (.A1(n_0_53), .A2(n_0_47), .A3(n_0_59), .ZN(n_0_111));
   NAND3_X1 i_0_126 (.A1(n_0_53), .A2(n_0_47), .A3(n_0_59), .ZN(n_0_112));
   NAND2_X1 i_0_152 (.A1(n_0_40), .A2(m[8]), .ZN(n_0_113));
   NAND2_X1 i_0_173 (.A1(n_0_112), .A2(n_0_113), .ZN(n_0_114));
   INV_X1 i_0_174 (.A(n_0_60), .ZN(n_0_115));
   NAND3_X1 i_0_177 (.A1(n_0_115), .A2(n_0_112), .A3(n_0_113), .ZN(n_0_116));
   INV_X1 i_0_179 (.A(n_0_116), .ZN(n_62));
   NAND2_X1 i_0_3 (.A1(n_0_126), .A2(r[0]), .ZN(n_0_117));
   INV_X1 i_0_21 (.A(n_0_117), .ZN(n_63));
   INV_X1 i_0_30 (.A(m[1]), .ZN(n_0_63));
   INV_X1 i_0_32 (.A(m[3]), .ZN(n_0_64));
   INV_X1 i_0_33 (.A(m[2]), .ZN(n_0_72));
   INV_X1 i_0_63 (.A(m[0]), .ZN(n_0_17));
   INV_X1 i_0_80 (.A(m[2]), .ZN(n_0_73));
   INV_X1 i_0_136 (.A(m[1]), .ZN(n_0_99));
   INV_X1 i_0_188 (.A(n_0_76), .ZN(n_0_127));
   INV_X1 i_0_189 (.A(n_0_136), .ZN(n_0_128));
   NAND2_X1 i_0_190 (.A1(n_0_127), .A2(n_0_128), .ZN(n_0_129));
   NAND3_X1 i_0_97 (.A1(n_0_163), .A2(n_0_129), .A3(r[0]), .ZN(n_0_131));
   INV_X1 i_0_185 (.A(n_0_131), .ZN(n_64));
   NAND3_X1 i_0_153 (.A1(n_0_167), .A2(n_0_168), .A3(n_0_169), .ZN(n_0_132));
   OAI21_X1 i_0_23 (.A(m[2]), .B1(m[0]), .B2(m[1]), .ZN(n_0_133));
   OAI21_X1 i_0_24 (.A(m[2]), .B1(m[0]), .B2(m[1]), .ZN(n_0_79));
   NAND4_X1 i_0_58 (.A1(n_0_106), .A2(n_0_67), .A3(n_0_68), .A4(n_0_66), 
      .ZN(n_0_139));
   NAND3_X1 i_0_59 (.A1(n_0_156), .A2(n_0_65), .A3(n_0_158), .ZN(n_0_140));
   INV_X1 i_0_154 (.A(m[3]), .ZN(n_0_100));
   NAND3_X1 i_0_94 (.A1(n_0_28), .A2(n_0_186), .A3(n_0_185), .ZN(n_0_80));
   INV_X1 i_0_41 (.A(m[0]), .ZN(n_0_148));
   INV_X1 i_0_43 (.A(m[1]), .ZN(n_0_149));
   INV_X1 i_0_62 (.A(m[2]), .ZN(n_0_150));
   NAND3_X1 i_0_77 (.A1(n_0_148), .A2(n_0_149), .A3(n_0_150), .ZN(n_0_151));
   INV_X1 i_0_88 (.A(m[3]), .ZN(n_0_152));
   NAND2_X1 i_0_112 (.A1(n_0_151), .A2(n_0_152), .ZN(n_0_153));
   NAND2_X1 i_0_144 (.A1(n_0_187), .A2(n_0_153), .ZN(n_65));
   NAND3_X1 i_0_61 (.A1(n_0_106), .A2(n_0_99), .A3(n_0_73), .ZN(n_0_155));
   NAND2_X1 i_0_66 (.A1(n_0_155), .A2(m[5]), .ZN(n_0_82));
   NAND2_X1 i_0_192 (.A1(n_0_20), .A2(n_0_24), .ZN(n_0_157));
   INV_X1 i_0_105 (.A(n_0_157), .ZN(n_0_90));
   INV_X1 i_0_42 (.A(n_0_93), .ZN(n_0_4));
   INV_X1 i_0_91 (.A(m[0]), .ZN(n_0_167));
   INV_X1 i_0_35 (.A(m[1]), .ZN(n_0_168));
   INV_X1 i_0_145 (.A(m[2]), .ZN(n_0_169));
   INV_X1 i_0_31 (.A(m[0]), .ZN(n_0_170));
   INV_X1 i_0_37 (.A(m[1]), .ZN(n_0_171));
   INV_X1 i_0_38 (.A(m[2]), .ZN(n_0_172));
   NAND3_X1 i_0_48 (.A1(n_0_170), .A2(n_0_171), .A3(n_0_172), .ZN(n_0_91));
   NAND3_X1 i_0_65 (.A1(n_0_25), .A2(n_0_98), .A3(n_0_138), .ZN(n_0_6));
   OAI21_X1 i_0_69 (.A(m[7]), .B1(n_0_140), .B2(n_0_139), .ZN(n_0_175));
   NAND2_X1 i_0_68 (.A1(n_0_100), .A2(n_0_17), .ZN(n_0_179));
   NAND2_X1 i_0_85 (.A1(n_0_179), .A2(m[5]), .ZN(n_0_95));
   NAND4_X1 i_0_64 (.A1(n_0_26), .A2(n_0_22), .A3(n_0_41), .A4(n_0_15), .ZN(
      n_0_70));
   INV_X1 i_0_92 (.A(n_0_70), .ZN(n_0_16));
   INV_X1 i_0_195 (.A(m[10]), .ZN(n_0_45));
   INV_X1 i_0_197 (.A(m[9]), .ZN(n_0_94));
   INV_X1 i_0_209 (.A(m[8]), .ZN(n_0_103));
   INV_X1 i_0_210 (.A(m[11]), .ZN(n_0_104));
   NOR2_X1 i_0_98 (.A1(m[0]), .A2(m[1]), .ZN(n_0_165));
   NOR2_X1 i_0_101 (.A1(m[5]), .A2(m[3]), .ZN(n_0_166));
   NOR2_X1 i_0_103 (.A1(m[2]), .A2(m[4]), .ZN(n_0_181));
   NAND3_X1 i_0_109 (.A1(n_0_165), .A2(n_0_166), .A3(n_0_181), .ZN(n_0_96));
   NAND4_X1 i_0_54 (.A1(n_0_65), .A2(n_0_67), .A3(n_0_68), .A4(n_0_66), .ZN(
      n_0_30));
   INV_X1 i_0_198 (.A(m[1]), .ZN(n_0_81));
   INV_X1 i_0_164 (.A(m[1]), .ZN(n_0_186));
   NAND3_X1 i_0_184 (.A1(n_0_197), .A2(n_0_198), .A3(n_0_90), .ZN(n_0_159));
   NAND4_X1 i_0_175 (.A1(n_0_143), .A2(n_0_144), .A3(n_0_145), .A4(n_0_146), 
      .ZN(n_0_102));
   NAND2_X1 i_0_180 (.A1(n_0_102), .A2(m[4]), .ZN(n_0_105));
   NAND3_X1 i_0_106 (.A1(n_0_197), .A2(n_0_198), .A3(n_0_90), .ZN(n_0_118));
   INV_X1 i_0_108 (.A(n_0_118), .ZN(n_0_122));
   INV_X1 i_0_123 (.A(n_0_48), .ZN(n_66));
   NAND3_X1 i_0_125 (.A1(n_0_82), .A2(n_0_95), .A3(n_0_96), .ZN(n_0_48));
   NAND4_X1 i_0_159 (.A1(n_0_82), .A2(n_0_95), .A3(r[0]), .A4(n_0_96), .ZN(
      n_0_124));
   INV_X1 i_0_204 (.A(n_0_124), .ZN(n_67));
   NAND4_X1 i_0_100 (.A1(n_0_143), .A2(n_0_144), .A3(n_0_145), .A4(n_0_146), 
      .ZN(n_0_76));
   NAND3_X1 i_0_113 (.A1(n_0_156), .A2(n_0_158), .A3(n_0_106), .ZN(n_0_136));
   NAND3_X1 i_0_115 (.A1(n_0_23), .A2(n_0_27), .A3(n_0_73), .ZN(n_0_161));
   NAND3_X1 i_0_120 (.A1(n_0_61), .A2(n_0_44), .A3(n_0_62), .ZN(n_0_162));
   INV_X1 i_0_121 (.A(m[0]), .ZN(n_0_143));
   INV_X1 i_0_122 (.A(m[1]), .ZN(n_0_144));
   INV_X1 i_0_138 (.A(m[3]), .ZN(n_0_145));
   INV_X1 i_0_140 (.A(m[2]), .ZN(n_0_146));
   INV_X1 i_0_141 (.A(m[6]), .ZN(n_0_156));
   INV_X1 i_0_143 (.A(m[5]), .ZN(n_0_158));
   INV_X1 i_0_181 (.A(m[4]), .ZN(n_0_106));
   NAND3_X1 i_0_163 (.A1(n_0_23), .A2(n_0_61), .A3(n_0_73), .ZN(n_0_109));
   NAND3_X1 i_0_178 (.A1(n_0_27), .A2(n_0_62), .A3(n_0_44), .ZN(n_0_119));
   NOR2_X1 i_0_219 (.A1(m[0]), .A2(m[1]), .ZN(n_0_120));
   NOR2_X1 i_0_220 (.A1(m[5]), .A2(m[3]), .ZN(n_0_123));
   NOR2_X1 i_0_221 (.A1(m[2]), .A2(m[4]), .ZN(n_0_154));
   NAND3_X1 i_0_99 (.A1(n_0_22), .A2(n_0_63), .A3(n_0_15), .ZN(n_0_19));
   INV_X1 i_0_111 (.A(n_0_19), .ZN(n_0_25));
   INV_X1 i_0_176 (.A(m[6]), .ZN(n_0_160));
   NAND4_X1 i_0_217 (.A1(n_0_120), .A2(n_0_123), .A3(n_0_154), .A4(n_0_160), 
      .ZN(n_0_173));
   INV_X1 i_0_218 (.A(n_0_109), .ZN(n_0_180));
   INV_X1 i_0_222 (.A(n_0_119), .ZN(n_0_182));
   NAND3_X1 i_0_223 (.A1(n_0_173), .A2(n_0_180), .A3(n_0_182), .ZN(n_0_184));
   NAND3_X1 i_0_224 (.A1(n_0_120), .A2(n_0_123), .A3(n_0_154), .ZN(n_0_188));
   NAND2_X1 i_0_225 (.A1(n_0_188), .A2(n_0_160), .ZN(n_0_189));
   NAND2_X1 i_0_226 (.A1(n_0_184), .A2(n_0_189), .ZN(n_68));
   NAND3_X1 i_0_127 (.A1(n_0_64), .A2(n_0_72), .A3(n_0_41), .ZN(n_0_134));
   INV_X1 i_0_135 (.A(n_0_134), .ZN(n_0_138));
   INV_X1 i_0_10 (.A(n_0_177), .ZN(n_69));
   NAND2_X1 i_0_15 (.A1(n_0_6), .A2(n_0_175), .ZN(n_0_177));
   NAND3_X1 i_0_84 (.A1(n_0_6), .A2(n_0_175), .A3(r[0]), .ZN(n_0_176));
   INV_X1 i_0_93 (.A(n_0_176), .ZN(n_70));
   INV_X1 i_0_211 (.A(n_0_110), .ZN(n_71));
   INV_X1 i_0_90 (.A(m[2]), .ZN(n_0_174));
   INV_X1 i_0_124 (.A(m[2]), .ZN(n_0_185));
   NAND4_X1 i_0_199 (.A1(n_0_28), .A2(n_0_81), .A3(m[3]), .A4(n_0_174), .ZN(
      n_0_187));
   OAI21_X1 i_0_83 (.A(m[6]), .B1(n_0_161), .B2(n_0_162), .ZN(n_0_163));
   NAND3_X1 i_0_67 (.A1(n_0_76), .A2(r[0]), .A3(n_0_75), .ZN(n_0_135));
   INV_X1 i_0_82 (.A(n_0_135), .ZN(n_72));
   NAND2_X1 i_0_51 (.A1(n_0_91), .A2(n_0_79), .ZN(n_0_125));
   INV_X1 i_0_56 (.A(n_0_125), .ZN(n_0_126));
   NAND3_X1 i_0_118 (.A1(n_0_192), .A2(n_0_197), .A3(n_0_198), .ZN(n_0_71));
   INV_X1 i_0_119 (.A(m[11]), .ZN(n_0_92));
   INV_X1 i_0_201 (.A(n_0_192), .ZN(n_0_101));
   INV_X1 i_0_207 (.A(n_0_92), .ZN(n_0_137));
   INV_X1 i_0_206 (.A(m[10]), .ZN(n_0_147));
   INV_X1 i_0_208 (.A(m[9]), .ZN(n_0_164));
   INV_X1 i_0_213 (.A(m[8]), .ZN(n_0_183));
   NAND3_X1 i_0_214 (.A1(n_0_147), .A2(n_0_164), .A3(n_0_183), .ZN(n_0_191));
   INV_X1 i_0_227 (.A(n_0_191), .ZN(n_0_192));
   NAND3_X1 i_0_166 (.A1(n_0_16), .A2(n_0_4), .A3(n_0_69), .ZN(n_0_194));
   NAND2_X1 i_0_182 (.A1(n_0_101), .A2(m[11]), .ZN(n_0_195));
   NAND3_X1 i_0_183 (.A1(n_0_199), .A2(n_0_194), .A3(n_0_195), .ZN(n_0_10));
   INV_X1 i_0_155 (.A(n_0_30), .ZN(n_0_197));
   INV_X1 i_0_193 (.A(n_0_0), .ZN(n_0_198));
   OAI21_X1 i_0_194 (.A(n_0_137), .B1(n_0_30), .B2(n_0_0), .ZN(n_0_199));
   INV_X1 i_0_71 (.A(n_0_7), .ZN(n_73));
   INV_X1 i_0_75 (.A(r[0]), .ZN(n_0_54));
   NOR2_X1 i_0_78 (.A1(n_0_7), .A2(n_0_54), .ZN(n_74));
   NAND3_X1 i_0_215 (.A1(n_0_215), .A2(n_0_105), .A3(r[0]), .ZN(n_0_110));
   NAND2_X1 i_0_216 (.A1(n_0_107), .A2(n_0_121), .ZN(n_0_130));
   NAND4_X1 i_0_202 (.A1(n_0_45), .A2(n_0_104), .A3(n_0_103), .A4(n_0_94), 
      .ZN(n_0_141));
   INV_X1 i_0_203 (.A(n_0_141), .ZN(n_0_69));
   INV_X1 i_0_81 (.A(n_0_193), .ZN(n_0_201));
   NAND3_X1 i_0_187 (.A1(n_0_16), .A2(n_0_4), .A3(n_0_69), .ZN(n_0_193));
   INV_X1 i_0_200 (.A(n_0_4), .ZN(n_0_202));
   INV_X1 i_0_229 (.A(m[12]), .ZN(n_0_203));
   NAND3_X1 i_0_230 (.A1(n_0_202), .A2(n_0_16), .A3(n_0_203), .ZN(n_0_204));
   INV_X1 i_0_231 (.A(n_0_16), .ZN(n_0_205));
   NAND2_X1 i_0_232 (.A1(n_0_205), .A2(n_0_203), .ZN(n_0_206));
   NAND2_X1 i_0_233 (.A1(n_0_204), .A2(n_0_206), .ZN(n_0_207));
   INV_X1 i_0_234 (.A(n_0_207), .ZN(n_0_208));
   XNOR2_X1 i_0_235 (.A(n_0_69), .B(n_0_203), .ZN(n_0_209));
   NAND2_X1 i_0_236 (.A1(n_0_16), .A2(n_0_4), .ZN(n_0_210));
   OAI21_X1 i_0_237 (.A(n_0_208), .B1(n_0_209), .B2(n_0_210), .ZN(n_75));
   INV_X1 i_0_205 (.A(n_0_9), .ZN(n_0_78));
   NOR2_X1 i_0_228 (.A1(m[12]), .A2(m[13]), .ZN(n_0_83));
   NAND2_X1 i_0_238 (.A1(n_0_78), .A2(n_0_83), .ZN(n_0_196));
   INV_X1 i_0_102 (.A(n_0_10), .ZN(n_76));
   INV_X1 i_0_161 (.A(n_0_10), .ZN(n_0_200));
   NAND2_X1 i_0_186 (.A1(n_0_200), .A2(n_0_3), .ZN(n_0_211));
   INV_X1 i_0_239 (.A(n_0_211), .ZN(n_77));
   INV_X1 i_0_57 (.A(n_0_178), .ZN(n_0_107));
   INV_X1 i_0_165 (.A(n_0_190), .ZN(n_0_121));
   NAND2_X1 i_0_191 (.A1(n_0_100), .A2(n_0_17), .ZN(n_0_178));
   NAND3_X1 i_0_196 (.A1(n_0_99), .A2(n_0_73), .A3(n_0_106), .ZN(n_0_190));
   NAND3_X1 i_0_212 (.A1(n_0_99), .A2(n_0_106), .A3(n_0_100), .ZN(n_0_142));
   INV_X1 i_0_240 (.A(n_0_142), .ZN(n_0_212));
   NAND2_X1 i_0_241 (.A1(n_0_17), .A2(n_0_73), .ZN(n_0_213));
   INV_X1 i_0_242 (.A(n_0_213), .ZN(n_0_214));
   NAND2_X1 i_0_243 (.A1(n_0_212), .A2(n_0_214), .ZN(n_0_215));
   NAND2_X1 i_5_0 (.A1(n_5_4727), .A2(n_5_45), .ZN(n_5_0));
   INV_X1 i_5_1 (.A(n_5_0), .ZN(n_5_1));
   AOI21_X1 i_5_2 (.A(n_5_1), .B1(n_5_4591), .B2(n_5_15), .ZN(n_5_2));
   INV_X1 i_5_3 (.A(n_5_4606), .ZN(n_5_3));
   INV_X1 i_5_4 (.A(r[10]), .ZN(n_5_4));
   NAND2_X1 i_5_5 (.A1(n_5_4), .A2(r[9]), .ZN(n_5_5));
   OAI21_X1 i_5_6 (.A(n_5_2), .B1(n_5_3), .B2(n_5_5), .ZN(n_78));
   NAND2_X1 i_5_7 (.A1(n_5_4592), .A2(n_5_15), .ZN(n_5_6));
   NAND2_X1 i_5_8 (.A1(n_5_4670), .A2(n_5_14), .ZN(n_5_7));
   NAND2_X1 i_5_9 (.A1(n_5_130), .A2(n_5_45), .ZN(n_5_8));
   NAND3_X1 i_5_10 (.A1(n_5_6), .A2(n_5_7), .A3(n_5_8), .ZN(n_79));
   NAND2_X1 i_5_11 (.A1(n_5_4593), .A2(n_5_15), .ZN(n_5_9));
   NAND2_X1 i_5_12 (.A1(n_5_4807), .A2(n_5_14), .ZN(n_5_10));
   NAND2_X1 i_5_13 (.A1(n_5_4610), .A2(n_5_45), .ZN(n_5_11));
   NAND3_X1 i_5_14 (.A1(n_5_9), .A2(n_5_10), .A3(n_5_11), .ZN(n_80));
   NAND2_X1 i_5_17 (.A1(n_5_4345), .A2(n_5_45), .ZN(n_5_13));
   NAND2_X1 i_5_21 (.A1(n_5_4307), .A2(n_5_45), .ZN(n_5_17));
   NAND3_X1 i_5_22 (.A1(n_5_4344), .A2(n_5_4616), .A3(n_5_17), .ZN(n_81));
   NAND2_X1 i_5_15 (.A1(n_5_4595), .A2(n_5_15), .ZN(n_5_18));
   NAND2_X1 i_5_19 (.A1(n_5_4607), .A2(n_5_14), .ZN(n_5_19));
   NAND2_X1 i_5_25 (.A1(n_5_4679), .A2(n_5_45), .ZN(n_5_20));
   NAND3_X1 i_5_23 (.A1(n_5_18), .A2(n_5_19), .A3(n_5_20), .ZN(n_82));
   NAND2_X1 i_5_26 (.A1(n_5_4596), .A2(n_5_15), .ZN(n_5_21));
   NAND2_X1 i_5_29 (.A1(n_5_711), .A2(n_5_45), .ZN(n_5_23));
   NAND3_X1 i_5_27 (.A1(n_5_21), .A2(n_5_4756), .A3(n_5_23), .ZN(n_83));
   NAND2_X1 i_5_33 (.A1(n_5_3961), .A2(n_5_45), .ZN(n_5_22));
   NAND2_X1 i_5_30 (.A1(n_5_4523), .A2(n_5_45), .ZN(n_5_24));
   NAND2_X1 i_5_39 (.A1(n_5_4598), .A2(n_5_15), .ZN(n_5_30));
   NAND2_X1 i_5_16 (.A1(n_5_4611), .A2(n_5_14), .ZN(n_5_31));
   NAND2_X1 i_5_41 (.A1(n_5_3856), .A2(n_5_45), .ZN(n_5_32));
   NAND3_X1 i_5_42 (.A1(n_5_30), .A2(n_5_31), .A3(n_5_32), .ZN(n_84));
   NAND2_X1 i_5_20 (.A1(n_5_4772), .A2(n_5_15), .ZN(n_5_33));
   NAND2_X1 i_5_28 (.A1(n_5_4612), .A2(n_5_14), .ZN(n_5_34));
   NAND2_X1 i_5_45 (.A1(n_5_4509), .A2(n_5_45), .ZN(n_5_35));
   NAND3_X1 i_5_31 (.A1(n_5_33), .A2(n_5_34), .A3(n_5_35), .ZN(n_85));
   NAND2_X1 i_5_49 (.A1(n_5_4635), .A2(n_5_45), .ZN(n_5_25));
   INV_X1 i_5_51 (.A(r[9]), .ZN(n_5_39));
   NOR2_X1 i_5_52 (.A1(r[10]), .A2(n_5_39), .ZN(n_5_14));
   NAND2_X1 i_5_53 (.A1(n_5_4614), .A2(n_5_14), .ZN(n_5_41));
   NAND2_X1 i_5_54 (.A1(r[10]), .A2(n_5_39), .ZN(n_5_42));
   INV_X1 i_5_55 (.A(n_5_42), .ZN(n_5_15));
   NAND2_X1 i_5_56 (.A1(n_5_4601), .A2(n_5_15), .ZN(n_5_44));
   XNOR2_X1 i_5_57 (.A(r[10]), .B(r[9]), .ZN(n_5_45));
   NAND2_X1 i_5_58 (.A1(n_5_4672), .A2(n_5_45), .ZN(n_5_46));
   NAND3_X1 i_5_59 (.A1(n_5_41), .A2(n_5_44), .A3(n_5_46), .ZN(n_86));
   BUF_X1 rt_shieldBuf__2__2__19 (.A(n_5_4727), .Z(n_5_12));
   XOR2_X1 i_5_60 (.A(m[0]), .B(n_5_12), .Z(n_5_4591));
   XOR2_X1 i_5_61 (.A(n_5_98), .B(n_5_40), .Z(n_5_4592));
   NAND2_X1 i_5_62 (.A1(n_5_139), .A2(n_5_97), .ZN(n_5_40));
   XNOR2_X1 i_5_40 (.A(n_5_121), .B(n_5_138), .ZN(n_5_4593));
   OAI21_X1 i_5_36 (.A(n_5_47), .B1(n_5_120), .B2(n_5_58), .ZN(n_5_16));
   OAI21_X1 i_5_64 (.A(n_5_152), .B1(n_5_151), .B2(n_5_58), .ZN(n_5_47));
   XOR2_X1 i_5_24 (.A(n_5_142), .B(n_5_48), .Z(n_5_4595));
   NAND2_X1 i_5_35 (.A1(n_5_4675), .A2(n_5_4676), .ZN(n_5_48));
   XOR2_X1 i_5_38 (.A(n_5_56), .B(n_5_4718), .Z(n_5_4596));
   XNOR2_X1 i_5_37 (.A(n_5_4552), .B(n_5_83), .ZN(n_5_27));
   XNOR2_X1 i_5_70 (.A(n_5_4734), .B(n_5_145), .ZN(n_5_4598));
   OAI21_X1 i_5_50 (.A(n_5_78), .B1(n_5_49), .B2(n_5_64), .ZN(n_5_37));
   NAND2_X1 i_5_66 (.A1(n_5_65), .A2(n_5_55), .ZN(n_5_49));
   NAND2_X1 i_5_75 (.A1(n_5_50), .A2(n_5_52), .ZN(n_5_4601));
   OAI21_X1 i_5_76 (.A(n_5_54), .B1(n_5_150), .B2(n_5_51), .ZN(n_5_50));
   NOR2_X1 i_5_77 (.A1(n_5_4672), .A2(n_75), .ZN(n_5_51));
   NAND3_X1 i_5_78 (.A1(n_5_67), .A2(n_5_148), .A3(n_5_53), .ZN(n_5_52));
   INV_X1 i_5_79 (.A(n_5_54), .ZN(n_5_53));
   AOI21_X1 i_5_80 (.A(n_5_64), .B1(n_5_55), .B2(n_5_65), .ZN(n_5_54));
   NAND2_X1 i_5_81 (.A1(n_5_63), .A2(n_5_115), .ZN(n_5_55));
   NAND2_X1 i_5_43 (.A1(n_5_57), .A2(n_5_4675), .ZN(n_5_56));
   NAND2_X1 i_5_44 (.A1(n_5_142), .A2(n_5_4676), .ZN(n_5_57));
   NOR2_X1 i_5_46 (.A1(n_5_4345), .A2(n_65), .ZN(n_5_58));
   INV_X1 i_5_47 (.A(n_5_85), .ZN(n_5_59));
   NAND2_X1 i_5_87 (.A1(n_5_68), .A2(n_5_69), .ZN(n_5_67));
   INV_X1 i_5_88 (.A(n_5_4672), .ZN(n_5_68));
   INV_X1 i_5_89 (.A(n_75), .ZN(n_5_69));
   NAND2_X1 i_5_73 (.A1(n_5_711), .A2(n_5_3185), .ZN(n_5_61));
   NOR2_X1 i_5_74 (.A1(n_5_711), .A2(n_5_3185), .ZN(n_5_62));
   NAND2_X1 i_5_84 (.A1(n_5_4773), .A2(n_5_116), .ZN(n_5_63));
   NOR2_X1 i_5_82 (.A1(n_5_4635), .A2(n_76), .ZN(n_5_64));
   NAND2_X1 i_5_86 (.A1(n_5_4635), .A2(n_76), .ZN(n_5_65));
   XNOR2_X1 i_5_83 (.A(n_5_4635), .B(n_76), .ZN(n_5_66));
   INV_X1 i_5_93 (.A(n_5_116), .ZN(n_5_70));
   INV_X1 i_5_98 (.A(n_5_4509), .ZN(n_5_71));
   INV_X1 i_5_99 (.A(n_73), .ZN(n_5_72));
   NAND2_X1 i_5_94 (.A1(n_5_71), .A2(n_5_72), .ZN(n_5_73));
   NAND2_X1 i_5_95 (.A1(n_5_70), .A2(n_5_73), .ZN(n_5_74));
   INV_X1 i_5_96 (.A(n_5_3706), .ZN(n_5_75));
   NAND2_X1 i_5_97 (.A1(n_5_73), .A2(n_5_75), .ZN(n_5_76));
   OAI21_X1 i_5_85 (.A(n_5_74), .B1(n_5_4724), .B2(n_5_76), .ZN(n_5_77));
   NAND2_X1 i_5_90 (.A1(n_5_66), .A2(n_5_77), .ZN(n_5_78));
   INV_X1 i_5_107 (.A(n_60), .ZN(n_5_80));
   OR2_X1 i_5_65 (.A1(n_5_4307), .A2(n_58), .ZN(n_5_84));
   NAND2_X1 i_5_48 (.A1(n_5_4307), .A2(n_58), .ZN(n_5_85));
   INV_X1 i_5_32 (.A(n_5_4551), .ZN(n_5_26));
   INV_X1 i_5_67 (.A(n_5_4541), .ZN(n_5_36));
   AOI21_X1 i_5_71 (.A(n_5_62), .B1(n_5_56), .B2(n_5_61), .ZN(n_5_83));
   NAND2_X1 i_5_100 (.A1(n_5_4381), .A2(n_5_80), .ZN(n_5_91));
   NAND2_X1 i_5_101 (.A1(n_5_4523), .A2(n_60), .ZN(n_5_92));
   AOI21_X1 i_5_102 (.A(n_5_62), .B1(n_5_56), .B2(n_5_61), .ZN(n_5_93));
   NAND2_X1 i_5_126 (.A1(n_5_130), .A2(n_5_4701), .ZN(n_5_97));
   NAND2_X1 i_5_127 (.A1(n_5_4727), .A2(m[0]), .ZN(n_5_98));
   NAND2_X1 i_5_130 (.A1(n_5_4701), .A2(m[0]), .ZN(n_5_101));
   INV_X1 i_5_131 (.A(n_5_101), .ZN(n_5_86));
   NAND2_X1 i_5_132 (.A1(n_59), .A2(m[0]), .ZN(n_5_103));
   INV_X1 i_5_133 (.A(n_5_103), .ZN(n_5_104));
   NAND2_X1 i_5_91 (.A1(n_5_4727), .A2(n_5_104), .ZN(n_5_105));
   INV_X1 i_5_63 (.A(n_5_105), .ZN(n_5_28));
   NAND2_X1 i_5_136 (.A1(n_5_4701), .A2(n_59), .ZN(n_5_107));
   INV_X1 i_5_137 (.A(n_5_107), .ZN(n_5_108));
   NAND2_X1 i_5_138 (.A1(n_59), .A2(m[0]), .ZN(n_5_109));
   INV_X1 i_5_139 (.A(n_5_109), .ZN(n_5_110));
   NAND2_X1 i_5_140 (.A1(n_5_4701), .A2(n_5_110), .ZN(n_5_111));
   INV_X1 i_5_141 (.A(n_5_111), .ZN(n_5_112));
   NAND2_X1 i_5_113 (.A1(n_5_92), .A2(n_5_91), .ZN(n_5_113));
   XNOR2_X1 i_5_117 (.A(n_5_114), .B(n_5_113), .ZN(n_5_29));
   NOR2_X1 i_5_118 (.A1(n_5_4551), .A2(n_5_4546), .ZN(n_5_114));
   OR2_X1 i_5_145 (.A1(n_5_4509), .A2(n_73), .ZN(n_5_115));
   NAND2_X1 i_5_146 (.A1(n_5_4509), .A2(n_73), .ZN(n_5_116));
   INV_X1 i_5_129 (.A(n_5_151), .ZN(n_5_118));
   INV_X1 i_5_142 (.A(n_5_152), .ZN(n_5_119));
   NAND2_X1 i_5_124 (.A1(n_5_118), .A2(n_5_119), .ZN(n_5_120));
   XNOR2_X1 i_5_104 (.A(n_5_4610), .B(n_59), .ZN(n_5_121));
   NOR2_X1 i_5_154 (.A1(n_5_4701), .A2(n_59), .ZN(n_5_124));
   NAND2_X1 i_5_125 (.A1(n_5_4735), .A2(n_5_124), .ZN(n_5_43));
   INV_X1 i_5_158 (.A(n_59), .ZN(n_5_128));
   NAND2_X1 i_5_69 (.A1(n_5_4735), .A2(n_5_128), .ZN(n_5_129));
   INV_X1 i_5_72 (.A(n_5_129), .ZN(n_5_60));
   INV_X1 i_5_106 (.A(n_5_130), .ZN(n_5_79));
   NAND2_X1 i_5_108 (.A1(n_5_4727), .A2(n_5_112), .ZN(n_5_133));
   INV_X1 i_5_164 (.A(n_5_108), .ZN(n_5_134));
   NAND2_X1 i_5_110 (.A1(n_5_133), .A2(n_5_134), .ZN(n_5_81));
   INV_X1 i_5_114 (.A(n_5_133), .ZN(n_5_82));
   NOR2_X1 i_5_167 (.A1(n_5_130), .A2(n_5_4701), .ZN(n_5_137));
   AOI21_X1 i_5_115 (.A(n_5_137), .B1(n_5_97), .B2(n_5_98), .ZN(n_5_138));
   INV_X1 i_5_169 (.A(n_5_140), .ZN(n_5_139));
   NOR2_X1 i_5_134 (.A1(n_5_130), .A2(n_5_4701), .ZN(n_5_140));
   NOR2_X1 i_5_122 (.A1(n_5_4491), .A2(n_5_58), .ZN(n_5_141));
   OAI21_X1 i_5_135 (.A(n_5_84), .B1(n_5_59), .B2(n_5_141), .ZN(n_5_142));
   NOR2_X1 i_5_148 (.A1(n_5_4491), .A2(n_5_58), .ZN(n_5_87));
   AOI21_X1 i_5_109 (.A(n_5_147), .B1(n_5_4624), .B2(n_5_4641), .ZN(n_5_145));
   INV_X1 i_5_92 (.A(n_5_3956), .ZN(n_5_88));
   NOR2_X1 i_5_166 (.A1(n_5_4523), .A2(n_60), .ZN(n_5_147));
   NAND2_X1 i_5_179 (.A1(n_5_4672), .A2(n_75), .ZN(n_5_148));
   NAND2_X1 i_5_180 (.A1(n_5_4672), .A2(n_75), .ZN(n_5_149));
   INV_X1 i_5_181 (.A(n_5_149), .ZN(n_5_150));
   INV_X1 i_5_143 (.A(n_5_153), .ZN(n_5_151));
   NAND2_X1 i_5_147 (.A1(n_5_154), .A2(n_5_155), .ZN(n_5_152));
   NAND2_X1 i_5_162 (.A1(n_5_4345), .A2(n_65), .ZN(n_5_153));
   NAND3_X1 i_5_175 (.A1(n_5_4617), .A2(n_5_4610), .A3(n_5_4609), .ZN(n_5_154));
   OAI22_X1 i_5_177 (.A1(n_5_28), .A2(n_5_81), .B1(n_5_130), .B2(n_5_82), 
      .ZN(n_5_155));
   NAND2_X1 i_5_151 (.A1(n_5_4345), .A2(n_65), .ZN(n_5_89));
   INV_X1 i_5_192 (.A(n_5_161), .ZN(n_5_4606));
   XNOR2_X1 i_5_193 (.A(n_5_507), .B(m[0]), .ZN(n_5_161));
   INV_X1 i_5_194 (.A(n_5_205), .ZN(n_5_3855));
   XOR2_X1 i_5_105 (.A(n_5_198), .B(n_5_195), .Z(n_5_4607));
   NAND2_X1 i_5_187 (.A1(n_5_3914), .A2(n_5_4291), .ZN(n_5_100));
   XNOR2_X1 i_5_68 (.A(n_5_3945), .B(n_5_200), .ZN(n_5_117));
   XNOR2_X1 i_5_18 (.A(n_5_4732), .B(n_5_4493), .ZN(n_5_4611));
   XOR2_X1 i_5_103 (.A(n_5_173), .B(n_5_4485), .Z(n_5_4612));
   XNOR2_X1 i_5_171 (.A(n_5_688), .B(n_5_172), .ZN(n_5_38));
   NAND2_X1 i_5_186 (.A1(n_5_164), .A2(n_5_167), .ZN(n_5_4614));
   OAI21_X1 i_5_189 (.A(n_5_661), .B1(n_5_165), .B2(n_5_166), .ZN(n_5_164));
   INV_X1 i_5_190 (.A(n_5_168), .ZN(n_5_165));
   NOR2_X1 i_5_191 (.A1(n_5_4672), .A2(n_5_169), .ZN(n_5_166));
   NAND3_X1 i_5_202 (.A1(n_5_170), .A2(n_5_659), .A3(n_5_168), .ZN(n_5_167));
   NAND2_X1 i_5_203 (.A1(n_5_4672), .A2(n_5_169), .ZN(n_5_168));
   INV_X1 i_5_210 (.A(m[12]), .ZN(n_5_169));
   NAND2_X1 i_5_206 (.A1(n_5_171), .A2(m[12]), .ZN(n_5_170));
   INV_X1 i_5_207 (.A(n_5_4672), .ZN(n_5_171));
   INV_X1 i_5_211 (.A(n_5_172), .ZN(n_5_437));
   OAI21_X1 i_5_178 (.A(n_5_190), .B1(n_5_191), .B2(n_5_173), .ZN(n_5_172));
   OAI21_X1 i_5_111 (.A(n_5_193), .B1(n_5_4493), .B2(n_5_179), .ZN(n_5_173));
   NAND2_X1 i_5_174 (.A1(n_5_198), .A2(n_5_4677), .ZN(n_5_122));
   NAND2_X1 i_5_153 (.A1(n_5_4727), .A2(m[0]), .ZN(n_5_90));
   NAND2_X1 i_5_155 (.A1(n_5_130), .A2(m[1]), .ZN(n_5_94));
   INV_X1 i_5_182 (.A(n_5_3978), .ZN(n_5_178));
   INV_X1 i_5_184 (.A(n_5_194), .ZN(n_5_179));
   NOR2_X1 i_5_213 (.A1(n_5_4635), .A2(m[11]), .ZN(n_5_450));
   NAND2_X1 i_5_226 (.A1(n_5_3961), .A2(m[7]), .ZN(n_5_96));
   INV_X1 i_5_229 (.A(m[11]), .ZN(n_5_468));
   INV_X1 i_5_231 (.A(m[6]), .ZN(n_5_125));
   INV_X1 i_5_123 (.A(n_5_3975), .ZN(n_5_186));
   OR2_X1 i_5_188 (.A1(n_5_4307), .A2(m[4]), .ZN(n_5_187));
   NAND2_X1 i_5_198 (.A1(n_5_4509), .A2(m[10]), .ZN(n_5_190));
   NOR2_X1 i_5_205 (.A1(n_5_4509), .A2(m[10]), .ZN(n_5_191));
   OR2_X1 i_5_212 (.A1(n_5_3856), .A2(m[9]), .ZN(n_5_193));
   NAND2_X1 i_5_172 (.A1(n_5_3856), .A2(m[9]), .ZN(n_5_194));
   NAND2_X1 i_5_112 (.A1(n_5_4678), .A2(n_5_4677), .ZN(n_5_195));
   OR2_X1 i_5_204 (.A1(n_5_4679), .A2(m[5]), .ZN(n_5_126));
   OR2_X1 i_5_157 (.A1(n_5_4610), .A2(m[2]), .ZN(n_5_99));
   XNOR2_X1 i_5_159 (.A(n_5_4610), .B(m[2]), .ZN(n_5_102));
   OAI21_X1 i_5_152 (.A(n_5_187), .B1(n_5_178), .B2(n_5_202), .ZN(n_5_198));
   AOI21_X1 i_5_163 (.A(n_5_186), .B1(n_5_4808), .B2(n_5_4372), .ZN(n_5_106));
   AOI21_X1 i_5_150 (.A(n_5_3858), .B1(n_5_96), .B2(n_5_3955), .ZN(n_5_200));
   AOI21_X1 i_5_161 (.A(n_5_186), .B1(n_5_4808), .B2(n_5_4372), .ZN(n_5_202));
   NOR2_X1 i_5_168 (.A1(n_5_130), .A2(m[1]), .ZN(n_5_123));
   NOR2_X1 i_5_259 (.A1(n_5_130), .A2(m[1]), .ZN(n_5_205));
   NAND2_X1 i_5_260 (.A1(n_5_558), .A2(n_5_95), .ZN(n_5_206));
   NAND2_X1 i_5_261 (.A1(n_5_491), .A2(n_5_188), .ZN(n_5_207));
   NAND2_X1 i_5_262 (.A1(n_5_4518), .A2(n_5_3866), .ZN(n_5_208));
   NAND3_X1 i_5_263 (.A1(n_5_206), .A2(n_5_207), .A3(n_5_208), .ZN(n_87));
   NAND2_X1 i_5_220 (.A1(n_5_499), .A2(n_5_188), .ZN(n_5_127));
   NAND2_X1 i_5_221 (.A1(n_5_559), .A2(n_5_95), .ZN(n_5_131));
   NAND2_X1 i_5_266 (.A1(n_5_696), .A2(n_5_3866), .ZN(n_5_143));
   NAND2_X1 i_5_170 (.A1(n_5_492), .A2(n_5_188), .ZN(n_5_212));
   NAND2_X1 i_5_173 (.A1(n_5_572), .A2(n_5_95), .ZN(n_5_213));
   NAND2_X1 i_5_270 (.A1(n_5_4436), .A2(n_5_3866), .ZN(n_5_214));
   NAND3_X1 i_5_185 (.A1(n_5_212), .A2(n_5_213), .A3(n_5_214), .ZN(n_5_130));
   NAND2_X1 i_5_264 (.A1(n_5_494), .A2(n_5_188), .ZN(n_5_144));
   NAND2_X1 i_5_236 (.A1(n_5_3968), .A2(n_5_3866), .ZN(n_5_146));
   NAND2_X1 i_5_248 (.A1(n_5_4682), .A2(n_5_3866), .ZN(n_5_180));
   NAND2_X1 i_5_119 (.A1(n_5_561), .A2(n_5_95), .ZN(n_5_4620));
   NAND2_X1 i_5_120 (.A1(n_5_502), .A2(n_5_188), .ZN(n_5_4621));
   NAND2_X1 i_5_278 (.A1(n_5_4501), .A2(n_5_3866), .ZN(n_5_4622));
   NAND2_X1 i_5_274 (.A1(n_5_3930), .A2(n_5_3866), .ZN(n_5_132));
   NAND2_X1 i_5_232 (.A1(n_5_4748), .A2(n_5_3866), .ZN(n_5_3863));
   NAND2_X1 i_5_241 (.A1(n_5_4338), .A2(n_5_3866), .ZN(n_5_136));
   NAND2_X1 i_5_237 (.A1(n_5_565), .A2(n_5_95), .ZN(n_5_220));
   NAND2_X1 i_5_238 (.A1(n_5_3964), .A2(n_5_3866), .ZN(n_5_222));
   INV_X1 i_5_288 (.A(r[8]), .ZN(n_5_223));
   NAND2_X1 i_5_289 (.A1(r[9]), .A2(n_5_223), .ZN(n_5_224));
   INV_X1 i_5_290 (.A(n_5_224), .ZN(n_5_95));
   NOR2_X1 i_5_291 (.A1(r[9]), .A2(n_5_223), .ZN(n_5_188));
   XNOR2_X1 i_5_292 (.A(r[9]), .B(r[8]), .ZN(n_5_3866));
   NAND2_X1 i_5_293 (.A1(n_5_4740), .A2(n_5_3866), .ZN(n_5_227));
   INV_X1 i_5_294 (.A(m[1]), .ZN(n_5_3867));
   NAND2_X1 i_5_265 (.A1(n_5_696), .A2(m[1]), .ZN(n_5_228));
   INV_X1 i_5_296 (.A(m[2]), .ZN(n_5_3868));
   INV_X1 i_5_297 (.A(m[3]), .ZN(n_5_229));
   NAND2_X1 i_5_298 (.A1(n_5_651), .A2(n_5_229), .ZN(n_5_3869));
   INV_X1 i_5_299 (.A(m[4]), .ZN(n_5_230));
   INV_X1 i_5_300 (.A(m[5]), .ZN(n_5_231));
   INV_X1 i_5_301 (.A(m[6]), .ZN(n_5_177));
   INV_X1 i_5_302 (.A(n_5_3930), .ZN(n_5_157));
   INV_X1 i_5_303 (.A(m[7]), .ZN(n_5_158));
   INV_X1 i_5_305 (.A(n_5_4660), .ZN(n_5_159));
   INV_X1 i_5_306 (.A(m[8]), .ZN(n_5_160));
   INV_X1 i_5_308 (.A(m[9]), .ZN(n_5_3877));
   INV_X1 i_5_310 (.A(m[10]), .ZN(n_5_3879));
   INV_X1 i_5_311 (.A(m[11]), .ZN(n_5_233));
   NAND2_X1 i_5_225 (.A1(n_5_4340), .A2(n_5_233), .ZN(n_5_3880));
   NAND2_X1 i_5_313 (.A1(n_5_4338), .A2(m[11]), .ZN(n_5_234));
   INV_X1 i_5_314 (.A(n_5_3964), .ZN(n_5_235));
   INV_X1 i_5_315 (.A(m[12]), .ZN(n_5_236));
   NAND2_X1 i_5_316 (.A1(n_5_235), .A2(n_5_236), .ZN(n_5_237));
   NAND2_X1 i_5_317 (.A1(n_5_3964), .A2(m[12]), .ZN(n_5_238));
   NAND2_X1 i_5_246 (.A1(n_5_3881), .A2(n_5_280), .ZN(n_5_135));
   NAND3_X1 i_5_320 (.A1(n_5_4531), .A2(n_5_485), .A3(n_5_228), .ZN(n_5_3881));
   AOI21_X1 i_5_321 (.A(n_5_4264), .B1(n_5_508), .B2(n_5_298), .ZN(n_5_3882));
   NOR2_X1 i_5_322 (.A1(n_5_508), .A2(n_5_4264), .ZN(n_5_3883));
   NAND2_X1 i_5_323 (.A1(n_5_3903), .A2(n_5_4262), .ZN(n_5_241));
   NAND2_X1 i_5_324 (.A1(n_5_271), .A2(n_5_619), .ZN(n_5_162));
   NAND3_X1 i_5_325 (.A1(n_5_4583), .A2(n_5_619), .A3(n_5_4264), .ZN(n_5_163));
   AOI21_X1 i_5_128 (.A(n_5_4253), .B1(n_5_260), .B2(n_5_264), .ZN(n_5_3886));
   NAND2_X1 i_5_327 (.A1(n_5_4577), .A2(n_5_4431), .ZN(n_5_3887));
   INV_X1 i_5_239 (.A(n_5_3880), .ZN(n_5_244));
   NAND2_X1 i_5_329 (.A1(n_5_4251), .A2(n_5_749), .ZN(n_5_245));
   INV_X1 i_5_330 (.A(n_5_245), .ZN(n_5_246));
   NAND2_X1 i_5_242 (.A1(n_5_539), .A2(n_5_246), .ZN(n_5_247));
   NOR2_X1 i_5_247 (.A1(n_5_244), .A2(n_5_247), .ZN(n_5_3888));
   INV_X1 i_5_243 (.A(n_5_234), .ZN(n_5_3889));
   NAND2_X1 i_5_334 (.A1(n_5_4251), .A2(n_5_295), .ZN(n_5_248));
   INV_X1 i_5_335 (.A(n_5_248), .ZN(n_5_175));
   INV_X1 i_5_337 (.A(n_5_264), .ZN(n_5_176));
   INV_X1 i_5_340 (.A(n_5_238), .ZN(n_5_253));
   OAI21_X1 i_5_341 (.A(n_5_237), .B1(n_5_532), .B2(n_5_253), .ZN(n_5_254));
   INV_X1 i_5_342 (.A(m[0]), .ZN(n_5_255));
   XNOR2_X1 i_5_343 (.A(n_5_257), .B(n_5_255), .ZN(n_5_491));
   XNOR2_X1 i_5_216 (.A(n_5_268), .B(n_5_675), .ZN(n_5_492));
   XNOR2_X1 i_5_282 (.A(n_5_4748), .B(m[9]), .ZN(n_5_189));
   BUF_X1 rt_shieldBuf__2__2__11 (.A(n_5_4518), .Z(n_5_257));
   INV_X1 i_5_349 (.A(m[1]), .ZN(n_5_511));
   NAND2_X1 i_5_350 (.A1(n_5_696), .A2(n_5_511), .ZN(n_5_258));
   AND3_X1 i_5_351 (.A1(n_5_690), .A2(n_5_4527), .A3(n_5_258), .ZN(n_5_259));
   NOR2_X1 i_5_352 (.A1(n_5_259), .A2(n_5_287), .ZN(n_5_499));
   OAI21_X1 i_5_219 (.A(n_5_749), .B1(n_5_295), .B2(n_5_4785), .ZN(n_5_260));
   NAND2_X1 i_5_144 (.A1(n_5_297), .A2(n_5_619), .ZN(n_5_262));
   NAND2_X1 i_5_223 (.A1(n_5_274), .A2(n_5_262), .ZN(n_5_3893));
   NAND2_X1 i_5_307 (.A1(n_5_4748), .A2(m[9]), .ZN(n_5_264));
   NAND2_X1 i_5_359 (.A1(n_5_4501), .A2(m[6]), .ZN(n_5_181));
   NAND2_X1 i_5_360 (.A1(n_5_4501), .A2(m[6]), .ZN(n_5_266));
   INV_X1 i_5_269 (.A(n_5_281), .ZN(n_5_267));
   OAI21_X1 i_5_233 (.A(n_5_284), .B1(n_5_228), .B2(n_5_267), .ZN(n_5_268));
   NAND2_X1 i_5_345 (.A1(n_5_4478), .A2(n_5_3869), .ZN(n_5_269));
   INV_X1 i_5_364 (.A(m[11]), .ZN(n_5_512));
   INV_X1 i_5_368 (.A(n_5_4404), .ZN(n_5_271));
   NAND2_X1 i_5_196 (.A1(n_5_266), .A2(n_5_4404), .ZN(n_5_272));
   NAND2_X1 i_5_208 (.A1(n_5_294), .A2(n_5_177), .ZN(n_5_273));
   NAND2_X1 i_5_209 (.A1(n_5_272), .A2(n_5_273), .ZN(n_5_274));
   INV_X1 i_5_372 (.A(m[6]), .ZN(n_5_275));
   XNOR2_X1 i_5_121 (.A(n_5_4501), .B(n_5_275), .ZN(n_5_276));
   XNOR2_X1 i_5_149 (.A(n_5_4314), .B(n_5_276), .ZN(n_5_502));
   INV_X1 i_5_375 (.A(m[13]), .ZN(n_5_277));
   XNOR2_X1 i_5_376 (.A(n_5_4740), .B(n_5_277), .ZN(n_5_278));
   XNOR2_X1 i_5_309 (.A(n_5_254), .B(n_5_278), .ZN(n_5_279));
   INV_X1 i_5_378 (.A(m[5]), .ZN(n_5_3898));
   NAND2_X1 i_5_380 (.A1(n_5_4448), .A2(n_5_3868), .ZN(n_5_280));
   NAND2_X1 i_5_304 (.A1(n_5_4526), .A2(n_5_3867), .ZN(n_5_281));
   NAND2_X1 i_5_319 (.A1(n_5_4526), .A2(n_5_3867), .ZN(n_5_282));
   INV_X1 i_5_344 (.A(n_5_4527), .ZN(n_5_283));
   NAND2_X1 i_5_358 (.A1(n_5_282), .A2(n_5_283), .ZN(n_5_284));
   AOI21_X1 i_5_385 (.A(n_5_4602), .B1(n_5_3869), .B2(n_5_4478), .ZN(n_5_182));
   NAND2_X1 i_5_386 (.A1(n_5_4518), .A2(m[0]), .ZN(n_5_286));
   AOI21_X1 i_5_387 (.A(n_5_286), .B1(n_5_690), .B2(n_5_258), .ZN(n_5_287));
   NOR2_X1 i_5_388 (.A1(n_5_231), .A2(n_5_230), .ZN(n_5_288));
   INV_X1 i_5_389 (.A(n_5_663), .ZN(n_5_289));
   INV_X1 i_5_390 (.A(n_5_231), .ZN(n_5_290));
   AOI21_X1 i_5_391 (.A(n_5_288), .B1(n_5_289), .B2(n_5_290), .ZN(n_5_232));
   NAND2_X1 i_5_392 (.A1(n_5_663), .A2(n_5_230), .ZN(n_5_292));
   INV_X1 i_5_393 (.A(n_5_292), .ZN(n_5_270));
   INV_X1 i_5_353 (.A(n_5_4577), .ZN(n_5_295));
   NAND2_X1 i_5_346 (.A1(n_5_159), .A2(n_5_160), .ZN(n_5_4626));
   NAND3_X1 i_5_355 (.A1(n_5_4583), .A2(n_5_241), .A3(n_5_4250), .ZN(n_5_296));
   INV_X1 i_5_251 (.A(n_5_296), .ZN(n_5_297));
   NAND2_X1 i_5_363 (.A1(n_5_663), .A2(n_5_230), .ZN(n_5_298));
   NAND2_X1 i_5_400 (.A1(n_5_663), .A2(n_5_230), .ZN(n_5_299));
   INV_X1 i_5_401 (.A(n_5_299), .ZN(n_5_3903));
   NAND2_X1 i_5_402 (.A1(n_5_4187), .A2(n_5_335), .ZN(n_5_300));
   INV_X1 i_5_403 (.A(n_5_300), .ZN(n_5_301));
   AOI21_X1 i_5_404 (.A(n_5_301), .B1(n_5_3976), .B2(n_5_197), .ZN(n_5_302));
   INV_X1 i_5_405 (.A(n_5_350), .ZN(n_5_303));
   INV_X1 i_5_406 (.A(r[8]), .ZN(n_5_304));
   NAND2_X1 i_5_407 (.A1(n_5_304), .A2(r[7]), .ZN(n_5_305));
   OAI21_X1 i_5_408 (.A(n_5_302), .B1(n_5_303), .B2(n_5_305), .ZN(n_88));
   NAND2_X1 i_5_409 (.A1(n_5_4159), .A2(n_5_335), .ZN(n_5_306));
   INV_X1 i_5_410 (.A(n_5_306), .ZN(n_5_307));
   AOI21_X1 i_5_411 (.A(n_5_307), .B1(n_5_351), .B2(n_5_218), .ZN(n_5_3904));
   INV_X1 i_5_412 (.A(n_5_3999), .ZN(n_5_3905));
   NAND2_X1 i_5_361 (.A1(n_5_4566), .A2(n_5_335), .ZN(n_5_517));
   NAND2_X1 i_5_245 (.A1(n_5_4311), .A2(n_5_335), .ZN(n_5_3906));
   NAND2_X1 i_5_415 (.A1(n_5_4461), .A2(n_5_335), .ZN(n_5_3907));
   NAND2_X1 i_5_416 (.A1(n_5_4476), .A2(n_5_335), .ZN(n_5_520));
   NAND2_X1 i_5_417 (.A1(n_5_4208), .A2(n_5_335), .ZN(n_5_4627));
   NAND2_X1 i_5_418 (.A1(n_5_4170), .A2(n_5_335), .ZN(n_5_3910));
   NAND2_X1 i_5_421 (.A1(n_5_4762), .A2(n_5_335), .ZN(n_5_183));
   NAND2_X1 i_5_422 (.A1(n_5_419), .A2(n_5_335), .ZN(n_5_184));
   NAND2_X1 i_5_228 (.A1(n_5_408), .A2(n_5_218), .ZN(n_5_185));
   NAND2_X1 i_5_424 (.A1(n_5_4507), .A2(n_5_335), .ZN(n_5_192));
   NAND2_X1 i_5_426 (.A1(n_5_4778), .A2(n_5_335), .ZN(n_5_196));
   NAND2_X1 i_5_428 (.A1(n_5_616), .A2(n_5_335), .ZN(n_5_3916));
   NAND2_X1 i_5_429 (.A1(n_5_4359), .A2(n_5_335), .ZN(n_5_324));
   INV_X1 i_5_430 (.A(n_5_324), .ZN(n_5_217));
   INV_X1 i_5_434 (.A(r[7]), .ZN(n_5_329));
   NOR2_X1 i_5_435 (.A1(r[8]), .A2(n_5_329), .ZN(n_5_218));
   NAND2_X1 i_5_436 (.A1(r[8]), .A2(n_5_329), .ZN(n_5_3918));
   INV_X1 i_5_437 (.A(n_5_3918), .ZN(n_5_197));
   XNOR2_X1 i_5_438 (.A(r[8]), .B(r[7]), .ZN(n_5_335));
   NAND2_X1 i_5_439 (.A1(n_5_381), .A2(n_5_335), .ZN(n_5_221));
   NAND2_X1 i_5_156 (.A1(n_5_3993), .A2(n_5_197), .ZN(n_5_3920));
   INV_X1 i_5_441 (.A(n_5_343), .ZN(n_5_350));
   XNOR2_X1 i_5_442 (.A(n_5_400), .B(m[0]), .ZN(n_5_343));
   XNOR2_X1 i_5_443 (.A(n_5_4159), .B(n_5_344), .ZN(n_5_351));
   NAND2_X1 i_5_444 (.A1(n_5_345), .A2(n_5_383), .ZN(n_5_344));
   INV_X1 i_5_445 (.A(n_5_384), .ZN(n_5_345));
   XNOR2_X1 i_5_382 (.A(n_5_658), .B(n_5_472), .ZN(n_5_545));
   XNOR2_X1 i_5_447 (.A(n_5_4460), .B(n_5_463), .ZN(n_5_3921));
   XOR2_X1 i_5_244 (.A(n_5_457), .B(n_5_401), .Z(n_5_4631));
   NAND2_X1 i_5_348 (.A1(n_5_454), .A2(n_5_361), .ZN(n_5_360));
   NAND2_X1 i_5_365 (.A1(n_5_4507), .A2(m[10]), .ZN(n_5_361));
   AOI21_X1 i_5_165 (.A(n_5_4328), .B1(n_5_251), .B2(n_5_649), .ZN(n_5_225));
   NAND2_X1 i_5_454 (.A1(n_5_369), .A2(n_5_370), .ZN(n_5_226));
   INV_X1 i_5_455 (.A(n_5_4359), .ZN(n_5_369));
   INV_X1 i_5_456 (.A(m[13]), .ZN(n_5_370));
   INV_X1 i_5_460 (.A(m[14]), .ZN(n_5_242));
   INV_X1 i_5_462 (.A(n_5_381), .ZN(n_5_243));
   OAI21_X1 i_5_312 (.A(n_5_250), .B1(n_5_4359), .B2(m[13]), .ZN(n_5_249));
   OAI21_X1 i_5_328 (.A(n_5_409), .B1(n_5_4632), .B2(n_5_379), .ZN(n_5_250));
   INV_X1 i_5_331 (.A(n_5_412), .ZN(n_5_379));
   INV_X1 i_5_466 (.A(m[10]), .ZN(n_5_251));
   NAND2_X1 i_5_272 (.A1(n_5_4170), .A2(m[7]), .ZN(n_5_459));
   NAND3_X1 i_5_257 (.A1(n_5_4187), .A2(m[1]), .A3(m[0]), .ZN(n_5_383));
   AOI21_X1 i_5_268 (.A(m[1]), .B1(n_5_4187), .B2(m[0]), .ZN(n_5_384));
   INV_X1 i_5_295 (.A(n_5_4159), .ZN(n_5_385));
   INV_X1 i_5_176 (.A(n_5_4760), .ZN(n_5_386));
   NOR2_X1 i_5_332 (.A1(n_5_616), .A2(m[12]), .ZN(n_5_4632));
   NAND2_X1 i_5_473 (.A1(n_5_4359), .A2(m[13]), .ZN(n_5_252));
   INV_X1 i_5_474 (.A(m[6]), .ZN(n_5_390));
   NAND2_X1 i_5_475 (.A1(n_5_4208), .A2(m[6]), .ZN(n_5_399));
   BUF_X1 rt_shieldBuf__2__2__12 (.A(n_5_4187), .Z(n_5_400));
   AOI21_X1 i_5_276 (.A(n_5_386), .B1(n_5_4759), .B2(n_5_430), .ZN(n_5_401));
   INV_X1 i_5_477 (.A(n_5_419), .ZN(n_5_402));
   INV_X1 i_5_478 (.A(m[9]), .ZN(n_5_403));
   INV_X1 i_5_479 (.A(n_5_458), .ZN(n_5_404));
   OAI21_X1 i_5_480 (.A(n_5_404), .B1(n_5_4208), .B2(m[6]), .ZN(n_5_405));
   NOR2_X1 i_5_279 (.A1(n_5_405), .A2(n_5_554), .ZN(n_5_406));
   OAI21_X1 i_5_280 (.A(n_5_406), .B1(n_5_4170), .B2(m[7]), .ZN(n_5_407));
   XNOR2_X1 i_5_396 (.A(n_5_360), .B(n_5_449), .ZN(n_5_408));
   NAND2_X1 i_5_333 (.A1(n_5_616), .A2(m[12]), .ZN(n_5_409));
   NAND2_X1 i_5_258 (.A1(n_5_616), .A2(m[12]), .ZN(n_5_411));
   OAI21_X1 i_5_336 (.A(n_5_4257), .B1(n_5_3807), .B2(n_5_4328), .ZN(n_5_412));
   OAI21_X1 i_5_273 (.A(n_5_4257), .B1(n_5_3807), .B2(n_5_4328), .ZN(n_5_414));
   NAND2_X1 i_5_283 (.A1(n_5_4632), .A2(n_5_414), .ZN(n_5_4633));
   XNOR2_X1 i_5_286 (.A(n_5_414), .B(n_5_411), .ZN(n_5_4634));
   XNOR2_X1 i_5_397 (.A(n_5_4208), .B(n_5_390), .ZN(n_5_422));
   NAND2_X1 i_5_399 (.A1(n_5_422), .A2(n_5_554), .ZN(n_5_549));
   INV_X1 i_5_497 (.A(n_5_390), .ZN(n_5_3927));
   XNOR2_X1 i_5_420 (.A(n_5_4204), .B(n_5_458), .ZN(n_5_550));
   NAND3_X1 i_5_339 (.A1(n_5_407), .A2(n_5_471), .A3(n_5_459), .ZN(n_5_428));
   XNOR2_X1 i_5_347 (.A(n_5_4758), .B(n_5_428), .ZN(n_5_261));
   NAND3_X1 i_5_183 (.A1(n_5_407), .A2(n_5_471), .A3(n_5_459), .ZN(n_5_430));
   NAND2_X1 i_5_502 (.A1(n_5_4311), .A2(m[3]), .ZN(n_5_199));
   NOR2_X1 i_5_503 (.A1(n_5_4311), .A2(m[3]), .ZN(n_5_433));
   OAI21_X1 i_5_195 (.A(n_5_399), .B1(n_5_4205), .B2(n_5_554), .ZN(n_5_3928));
   OAI21_X1 i_5_505 (.A(n_5_399), .B1(n_5_4205), .B2(n_5_554), .ZN(n_5_475));
   NAND2_X1 i_5_377 (.A1(n_5_249), .A2(n_5_252), .ZN(n_5_263));
   NAND2_X1 i_5_200 (.A1(n_5_402), .A2(n_5_403), .ZN(n_5_441));
   NAND2_X1 i_5_215 (.A1(n_5_402), .A2(n_5_403), .ZN(n_5_442));
   NAND3_X1 i_5_217 (.A1(n_5_430), .A2(n_5_441), .A3(n_5_4759), .ZN(n_5_156));
   NAND2_X1 i_5_240 (.A1(n_5_442), .A2(n_5_386), .ZN(n_5_174));
   NAND2_X1 i_5_252 (.A1(n_5_419), .A2(m[9]), .ZN(n_5_239));
   NAND3_X1 i_5_476 (.A1(n_5_441), .A2(n_5_430), .A3(n_5_4759), .ZN(n_5_446));
   NAND2_X1 i_5_501 (.A1(n_5_442), .A2(n_5_386), .ZN(n_5_447));
   NAND2_X1 i_5_509 (.A1(n_5_419), .A2(m[9]), .ZN(n_5_448));
   NAND3_X1 i_5_510 (.A1(n_5_446), .A2(n_5_447), .A3(n_5_448), .ZN(n_5_449));
   NAND2_X1 i_5_362 (.A1(n_5_4566), .A2(m[2]), .ZN(n_5_503));
   NAND2_X1 i_5_514 (.A1(n_5_649), .A2(n_5_251), .ZN(n_5_454));
   XNOR2_X1 i_5_284 (.A(n_5_419), .B(m[9]), .ZN(n_5_457));
   NOR2_X1 i_5_431 (.A1(n_5_4476), .A2(m[5]), .ZN(n_5_458));
   AOI21_X1 i_5_527 (.A(n_5_433), .B1(n_5_4814), .B2(n_5_199), .ZN(n_5_463));
   NAND2_X1 i_5_529 (.A1(n_5_256), .A2(n_5_433), .ZN(n_5_466));
   NAND2_X1 i_5_530 (.A1(n_5_4812), .A2(n_5_466), .ZN(n_5_467));
   OR2_X1 i_5_531 (.A1(n_5_4170), .A2(m[7]), .ZN(n_5_518));
   NAND2_X1 i_5_532 (.A1(n_5_4208), .A2(m[6]), .ZN(n_5_469));
   INV_X1 i_5_370 (.A(n_5_469), .ZN(n_5_470));
   OAI21_X1 i_5_373 (.A(n_5_470), .B1(n_5_4170), .B2(m[7]), .ZN(n_5_471));
   AOI21_X1 i_5_414 (.A(n_5_384), .B1(n_5_385), .B2(n_5_383), .ZN(n_5_472));
   INV_X1 i_5_384 (.A(n_5_384), .ZN(n_5_473));
   NAND2_X1 i_5_413 (.A1(n_5_385), .A2(n_5_383), .ZN(n_5_474));
   NAND2_X1 i_5_446 (.A1(n_5_473), .A2(n_5_474), .ZN(n_5_522));
   NOR2_X1 i_5_539 (.A1(n_5_467), .A2(n_5_4302), .ZN(n_5_3934));
   NAND2_X1 i_5_540 (.A1(n_5_4476), .A2(m[5]), .ZN(n_5_477));
   NAND2_X1 i_5_457 (.A1(n_5_467), .A2(n_5_477), .ZN(n_5_478));
   NAND2_X1 i_5_458 (.A1(n_5_477), .A2(n_5_4302), .ZN(n_5_479));
   NAND2_X1 i_5_463 (.A1(n_5_478), .A2(n_5_479), .ZN(n_5_554));
   NAND2_X1 i_5_281 (.A1(n_5_4507), .A2(m[10]), .ZN(n_5_496));
   NAND3_X1 i_5_545 (.A1(n_5_3973), .A2(n_5_3972), .A3(n_5_3906), .ZN(n_5_484));
   NAND2_X1 i_5_546 (.A1(n_5_484), .A2(m[2]), .ZN(n_5_485));
   BUF_X1 rt_shieldBuf__2__2__14 (.A(n_5_4727), .Z(n_5_507));
   NAND2_X1 i_5_549 (.A1(n_5_269), .A2(n_5_353), .ZN(n_5_308));
   XNOR2_X1 i_5_481 (.A(n_5_308), .B(n_5_668), .ZN(n_5_494));
   NAND2_X1 i_5_483 (.A1(n_5_269), .A2(n_5_353), .ZN(n_5_508));
   INV_X1 i_5_552 (.A(m[12]), .ZN(n_5_309));
   XNOR2_X1 i_5_440 (.A(n_5_4421), .B(n_5_309), .ZN(n_5_265));
   NAND2_X1 i_5_464 (.A1(n_5_4635), .A2(m[11]), .ZN(n_5_556));
   NAND3_X1 i_5_448 (.A1(n_5_220), .A2(n_5_4789), .A3(n_5_222), .ZN(n_5_4635));
   NAND3_X1 i_5_366 (.A1(n_5_4789), .A2(n_5_220), .A3(n_5_222), .ZN(n_5_557));
   NAND2_X1 i_5_557 (.A1(n_5_339), .A2(n_5_320), .ZN(n_5_311));
   INV_X1 i_5_558 (.A(m[0]), .ZN(n_5_312));
   XNOR2_X1 i_5_559 (.A(n_5_313), .B(n_5_312), .ZN(n_5_558));
   XNOR2_X1 i_5_560 (.A(n_5_693), .B(n_5_314), .ZN(n_5_559));
   BUF_X1 rt_shieldBuf__2__2__17 (.A(n_5_4518), .Z(n_5_313));
   INV_X1 i_5_561 (.A(n_5_4520), .ZN(n_5_314));
   INV_X1 i_5_562 (.A(n_5_2568), .ZN(n_5_315));
   AOI21_X1 i_5_255 (.A(n_5_424), .B1(n_5_397), .B2(n_5_354), .ZN(n_5_201));
   AOI21_X1 i_5_197 (.A(n_5_346), .B1(n_5_365), .B2(n_5_394), .ZN(n_5_317));
   XOR2_X1 i_5_199 (.A(n_5_4504), .B(n_5_317), .Z(n_5_561));
   NOR2_X1 i_5_254 (.A1(n_5_389), .A2(n_5_416), .ZN(n_5_562));
   XNOR2_X1 i_5_287 (.A(n_5_603), .B(n_5_4514), .ZN(n_5_563));
   NAND2_X1 i_5_515 (.A1(n_5_417), .A2(n_5_391), .ZN(n_5_564));
   INV_X1 i_5_570 (.A(n_5_423), .ZN(n_5_318));
   AOI21_X1 i_5_571 (.A(n_5_318), .B1(n_5_358), .B2(n_5_391), .ZN(n_5_3938));
   XNOR2_X1 i_5_491 (.A(n_5_608), .B(n_5_4283), .ZN(n_5_565));
   XNOR2_X1 i_5_492 (.A(n_5_4740), .B(n_61), .ZN(n_5_319));
   BUF_X1 i_5_574 (.A(n_5_382), .Z(n_5_320));
   NAND2_X1 i_5_493 (.A1(n_5_3964), .A2(n_75), .ZN(n_5_321));
   INV_X1 i_5_576 (.A(n_5_3944), .ZN(n_5_322));
   INV_X1 i_5_578 (.A(n_60), .ZN(n_5_328));
   INV_X1 i_5_579 (.A(n_66), .ZN(n_5_330));
   NOR2_X1 i_5_356 (.A1(n_5_4748), .A2(n_55), .ZN(n_5_3939));
   INV_X1 i_5_581 (.A(n_55), .ZN(n_5_331));
   NOR2_X1 i_5_582 (.A1(n_5_4501), .A2(n_5_3185), .ZN(n_5_332));
   INV_X1 i_5_585 (.A(n_5_330), .ZN(n_5_3940));
   INV_X1 i_5_587 (.A(n_5_315), .ZN(n_5_337));
   NAND2_X1 i_5_468 (.A1(n_5_696), .A2(n_5_337), .ZN(n_5_338));
   BUF_X1 i_5_589 (.A(n_5_340), .Z(n_5_339));
   NAND2_X1 i_5_590 (.A1(n_5_426), .A2(n_5_331), .ZN(n_5_340));
   NAND2_X1 i_5_494 (.A1(n_5_4289), .A2(n_5_321), .ZN(n_5_341));
   XNOR2_X1 i_5_506 (.A(n_5_319), .B(n_5_341), .ZN(n_5_568));
   INV_X1 i_5_593 (.A(n_58), .ZN(n_5_342));
   NAND2_X1 i_5_594 (.A1(n_5_4501), .A2(n_5_3185), .ZN(n_5_285));
   NAND2_X1 i_5_596 (.A1(n_5_4338), .A2(n_76), .ZN(n_5_3941));
   NAND2_X1 i_5_357 (.A1(n_5_4650), .A2(n_5_328), .ZN(n_5_3942));
   NAND2_X1 i_5_598 (.A1(n_5_4650), .A2(n_5_328), .ZN(n_5_348));
   OAI21_X1 i_5_599 (.A(n_5_3997), .B1(n_5_4008), .B2(n_5_4009), .ZN(n_5_349));
   NAND2_X1 i_5_600 (.A1(n_5_348), .A2(n_5_349), .ZN(n_5_352));
   NAND2_X1 i_5_519 (.A1(n_5_352), .A2(n_5_4254), .ZN(n_5_3943));
   NAND2_X1 i_5_516 (.A1(n_5_285), .A2(n_5_332), .ZN(n_5_310));
   OAI21_X1 i_5_605 (.A(n_5_3951), .B1(n_5_3939), .B2(n_5_334), .ZN(n_5_356));
   INV_X1 i_5_606 (.A(n_5_356), .ZN(n_5_357));
   OAI21_X1 i_5_607 (.A(n_5_357), .B1(n_5_311), .B2(n_5_322), .ZN(n_5_358));
   OAI21_X1 i_5_369 (.A(n_5_3997), .B1(n_5_4009), .B2(n_5_4008), .ZN(n_5_3944));
   NAND2_X1 i_5_610 (.A1(n_5_431), .A2(n_5_4226), .ZN(n_5_359));
   INV_X1 i_5_611 (.A(n_5_431), .ZN(n_5_362));
   OAI21_X1 i_5_612 (.A(n_5_359), .B1(n_5_427), .B2(n_5_362), .ZN(n_5_323));
   INV_X1 i_5_613 (.A(n_5_342), .ZN(n_5_366));
   OAI21_X1 i_5_614 (.A(n_5_664), .B1(n_5_3968), .B2(n_5_366), .ZN(n_5_571));
   OAI21_X1 i_5_518 (.A(n_5_338), .B1(n_5_694), .B2(n_5_4520), .ZN(n_5_368));
   XNOR2_X1 i_5_528 (.A(n_5_679), .B(n_5_368), .ZN(n_5_572));
   NOR3_X1 i_5_256 (.A1(n_5_642), .A2(n_5_4226), .A3(n_5_4343), .ZN(n_5_371));
   NOR2_X1 i_5_214 (.A1(n_5_4682), .A2(n_66), .ZN(n_5_346));
   INV_X1 i_5_619 (.A(n_65), .ZN(n_5_380));
   INV_X1 i_5_620 (.A(n_5_336), .ZN(n_5_382));
   NAND2_X1 i_5_224 (.A1(n_5_4682), .A2(n_66), .ZN(n_5_365));
   INV_X1 i_5_354 (.A(n_5_4401), .ZN(n_5_388));
   NOR3_X1 i_5_371 (.A1(n_5_4503), .A2(n_5_371), .A3(n_5_388), .ZN(n_5_389));
   INV_X1 i_5_624 (.A(n_65), .ZN(n_5_203));
   INV_X1 i_5_625 (.A(n_5_380), .ZN(n_5_209));
   INV_X1 i_5_626 (.A(n_5_315), .ZN(n_5_577));
   OR2_X1 i_5_584 (.A1(n_5_4665), .A2(n_73), .ZN(n_5_391));
   NAND2_X1 i_5_485 (.A1(n_5_525), .A2(n_5_4403), .ZN(n_5_325));
   XNOR2_X1 i_5_486 (.A(n_5_413), .B(n_5_4682), .ZN(n_5_326));
   INV_X1 i_5_630 (.A(n_5_3968), .ZN(n_5_392));
   NAND2_X1 i_5_227 (.A1(n_5_392), .A2(n_5_342), .ZN(n_5_393));
   OAI21_X1 i_5_234 (.A(n_5_393), .B1(n_5_427), .B2(n_5_435), .ZN(n_5_394));
   NOR2_X1 i_5_633 (.A1(n_5_696), .A2(n_5_2568), .ZN(n_5_395));
   OAI21_X1 i_5_267 (.A(n_5_338), .B1(n_5_4520), .B2(n_5_395), .ZN(n_5_396));
   INV_X1 i_5_318 (.A(n_5_396), .ZN(n_5_397));
   NAND2_X1 i_5_636 (.A1(n_5_415), .A2(n_5_694), .ZN(n_5_398));
   INV_X1 i_5_637 (.A(n_5_398), .ZN(n_5_327));
   NOR2_X1 i_5_638 (.A1(n_5_4338), .A2(n_76), .ZN(n_5_3948));
   INV_X1 i_5_639 (.A(n_76), .ZN(n_5_580));
   XNOR2_X1 i_5_629 (.A(n_5_666), .B(n_5_3940), .ZN(n_5_413));
   NAND2_X1 i_5_641 (.A1(n_5_696), .A2(n_5_577), .ZN(n_5_415));
   NOR2_X1 i_5_374 (.A1(n_5_4501), .A2(n_5_3185), .ZN(n_5_416));
   INV_X1 i_5_643 (.A(n_5_3185), .ZN(n_5_3949));
   OAI211_X1 i_5_602 (.A(n_5_4423), .B(n_5_3951), .C1(n_5_3939), .C2(n_5_4515), 
      .ZN(n_5_417));
   NAND2_X1 i_5_645 (.A1(n_5_4665), .A2(n_73), .ZN(n_5_423));
   NOR2_X1 i_5_383 (.A1(n_5_4436), .A2(n_59), .ZN(n_5_424));
   INV_X1 i_5_647 (.A(n_59), .ZN(n_5_3950));
   INV_X1 i_5_648 (.A(n_5_4520), .ZN(n_5_425));
   NAND2_X1 i_5_395 (.A1(n_5_4748), .A2(n_55), .ZN(n_5_3951));
   INV_X1 i_5_650 (.A(n_5_4748), .ZN(n_5_426));
   INV_X1 i_5_651 (.A(n_55), .ZN(n_5_3952));
   INV_X1 i_5_652 (.A(n_5_331), .ZN(n_5_3953));
   OAI21_X1 i_5_235 (.A(n_5_4524), .B1(n_5_2184), .B2(n_5_4290), .ZN(n_5_427));
   OAI21_X1 i_5_654 (.A(n_5_4524), .B1(n_5_2184), .B2(n_5_4290), .ZN(n_5_3954));
   NAND2_X1 i_5_655 (.A1(n_5_3968), .A2(n_58), .ZN(n_5_431));
   NAND2_X1 i_5_656 (.A1(n_5_3968), .A2(n_58), .ZN(n_5_434));
   INV_X1 i_5_249 (.A(n_5_434), .ZN(n_5_435));
   NAND2_X1 i_5_642 (.A1(n_5_425), .A2(n_59), .ZN(n_5_333));
   INV_X1 i_5_661 (.A(m[3]), .ZN(n_5_3957));
   INV_X1 i_5_662 (.A(m[2]), .ZN(n_5_590));
   XNOR2_X1 i_5_489 (.A(n_5_4294), .B(n_5_571), .ZN(n_5_591));
   NAND2_X1 i_5_469 (.A1(n_5_591), .A2(n_5_95), .ZN(n_5_210));
   NAND2_X1 i_5_495 (.A1(n_5_550), .A2(n_5_549), .ZN(n_5_4636));
   INV_X1 i_5_666 (.A(n_5_218), .ZN(n_5_594));
   AOI21_X1 i_5_496 (.A(n_5_594), .B1(n_5_549), .B2(n_5_554), .ZN(n_5_4637));
   NAND3_X1 i_5_423 (.A1(n_5_4689), .A2(n_5_4690), .A3(n_5_184), .ZN(n_5_597));
   NAND2_X1 i_5_381 (.A1(n_5_597), .A2(n_60), .ZN(n_5_334));
   NOR2_X1 i_5_670 (.A1(n_5_597), .A2(n_60), .ZN(n_5_336));
   XNOR2_X1 i_5_201 (.A(n_5_597), .B(m[8]), .ZN(n_5_529));
   XNOR2_X1 i_5_427 (.A(n_5_3982), .B(n_73), .ZN(n_5_603));
   XNOR2_X1 i_5_432 (.A(n_5_3982), .B(m[10]), .ZN(n_5_3963));
   INV_X1 i_5_508 (.A(n_5_4421), .ZN(n_5_3964));
   INV_X1 i_5_676 (.A(n_75), .ZN(n_5_607));
   XNOR2_X1 i_5_553 (.A(n_5_4421), .B(n_5_607), .ZN(n_5_608));
   NAND2_X1 i_5_470 (.A1(n_5_545), .A2(n_5_218), .ZN(n_5_609));
   NAND2_X1 i_5_490 (.A1(n_5_3977), .A2(n_5_197), .ZN(n_5_610));
   XNOR2_X1 i_5_379 (.A(n_5_4638), .B(n_69), .ZN(n_5_617));
   XNOR2_X1 i_5_394 (.A(n_5_4638), .B(m[7]), .ZN(n_5_3965));
   NAND2_X1 i_5_686 (.A1(n_5_188), .A2(m[2]), .ZN(n_5_627));
   INV_X1 i_5_687 (.A(n_5_627), .ZN(n_5_628));
   NAND2_X1 i_5_498 (.A1(n_5_4796), .A2(n_5_628), .ZN(n_5_629));
   NAND2_X1 i_5_689 (.A1(n_5_95), .A2(m[2]), .ZN(n_5_630));
   INV_X1 i_5_690 (.A(n_5_630), .ZN(n_5_631));
   NAND2_X1 i_5_533 (.A1(n_5_4040), .A2(n_5_631), .ZN(n_5_632));
   INV_X1 i_5_692 (.A(n_5_4408), .ZN(n_5_633));
   NAND2_X1 i_5_693 (.A1(n_5_633), .A2(m[2]), .ZN(n_5_634));
   NAND3_X1 i_5_535 (.A1(n_5_629), .A2(n_5_632), .A3(n_5_634), .ZN(n_5_211));
   XNOR2_X1 i_5_419 (.A(n_5_562), .B(n_5_617), .ZN(n_5_636));
   NAND2_X1 i_5_499 (.A1(n_5_636), .A2(n_5_95), .ZN(n_5_347));
   NOR2_X1 i_5_425 (.A1(n_5_4682), .A2(n_66), .ZN(n_5_642));
   NAND2_X1 i_5_504 (.A1(n_5_3873), .A2(m[3]), .ZN(n_5_353));
   INV_X1 i_5_702 (.A(n_5_3873), .ZN(n_5_651));
   INV_X1 i_5_615 (.A(n_5_4566), .ZN(n_5_655));
   INV_X1 i_5_704 (.A(m[2]), .ZN(n_5_656));
   INV_X1 i_5_705 (.A(n_5_590), .ZN(n_5_657));
   OAI22_X1 i_5_616 (.A1(n_5_655), .A2(n_5_656), .B1(n_5_4566), .B2(n_5_657), 
      .ZN(n_5_658));
   AOI21_X1 i_5_554 (.A(n_5_450), .B1(n_5_556), .B2(n_5_437), .ZN(n_5_659));
   AOI21_X1 i_5_708 (.A(n_5_450), .B1(n_5_437), .B2(n_5_556), .ZN(n_5_660));
   INV_X1 i_5_556 (.A(n_5_660), .ZN(n_5_661));
   NAND3_X1 i_5_640 (.A1(n_5_4332), .A2(n_5_4480), .A3(n_5_520), .ZN(n_5_662));
   INV_X1 i_5_521 (.A(n_5_662), .ZN(n_5_663));
   NAND2_X1 i_5_712 (.A1(n_5_662), .A2(n_58), .ZN(n_5_664));
   NAND2_X1 i_5_713 (.A1(n_5_662), .A2(n_58), .ZN(n_5_3967));
   NAND2_X1 i_5_710 (.A1(n_5_662), .A2(n_58), .ZN(n_5_666));
   XNOR2_X1 i_5_715 (.A(n_5_662), .B(m[4]), .ZN(n_5_668));
   NAND3_X1 i_5_523 (.A1(n_5_4332), .A2(n_5_4480), .A3(n_5_520), .ZN(n_5_3968));
   NAND3_X1 i_5_621 (.A1(n_5_4730), .A2(n_5_4495), .A3(n_5_3916), .ZN(n_5_670));
   XNOR2_X1 i_5_627 (.A(n_5_670), .B(n_5_580), .ZN(n_5_671));
   XNOR2_X1 i_5_631 (.A(n_5_670), .B(n_5_512), .ZN(n_5_3969));
   XNOR2_X1 i_5_536 (.A(n_5_4449), .B(m[2]), .ZN(n_5_675));
   NAND2_X1 i_5_563 (.A1(n_5_4436), .A2(n_59), .ZN(n_5_354));
   XNOR2_X1 i_5_537 (.A(n_5_4449), .B(n_59), .ZN(n_5_679));
   NAND2_X1 i_5_723 (.A1(n_5_577), .A2(n_59), .ZN(n_5_682));
   INV_X1 i_5_724 (.A(n_5_682), .ZN(n_5_683));
   NAND2_X1 i_5_703 (.A1(n_5_696), .A2(n_5_683), .ZN(n_5_355));
   INV_X1 i_5_573 (.A(n_5_557), .ZN(n_5_685));
   INV_X1 i_5_727 (.A(m[11]), .ZN(n_5_686));
   INV_X1 i_5_728 (.A(n_5_468), .ZN(n_5_687));
   OAI22_X1 i_5_618 (.A1(n_5_685), .A2(n_5_686), .B1(n_5_557), .B2(n_5_687), 
      .ZN(n_5_688));
   NAND3_X1 i_5_538 (.A1(n_5_609), .A2(n_5_610), .A3(n_5_517), .ZN(n_5_3970));
   OR2_X1 i_5_731 (.A1(n_5_3970), .A2(n_5_511), .ZN(n_5_690));
   XNOR2_X1 i_5_733 (.A(n_5_3970), .B(n_5_2568), .ZN(n_5_693));
   NOR2_X1 i_5_543 (.A1(n_5_3970), .A2(n_5_2568), .ZN(n_5_694));
   NAND2_X1 i_5_706 (.A1(n_5_696), .A2(n_5_577), .ZN(n_5_3971));
   NAND3_X1 i_5_551 (.A1(n_5_609), .A2(n_5_610), .A3(n_5_517), .ZN(n_5_696));
   NAND2_X1 i_5_449 (.A1(n_5_563), .A2(n_5_95), .ZN(n_5_4639));
   NAND2_X1 i_5_450 (.A1(n_5_4665), .A2(n_5_3866), .ZN(n_5_4640));
   NAND2_X1 i_5_743 (.A1(n_5_4804), .A2(n_5_197), .ZN(n_5_3972));
   NAND2_X1 i_5_588 (.A1(n_5_4811), .A2(n_5_218), .ZN(n_5_3973));
   XNOR2_X1 i_5_632 (.A(n_5_564), .B(n_5_671), .ZN(n_5_710));
   NAND2_X1 i_5_451 (.A1(n_5_710), .A2(n_5_95), .ZN(n_5_363));
   INV_X1 i_5_749 (.A(m[3]), .ZN(n_5_592));
   NAND2_X1 i_5_750 (.A1(n_5_146), .A2(n_5_592), .ZN(n_5_712));
   INV_X1 i_5_722 (.A(n_5_712), .ZN(n_5_713));
   NAND3_X1 i_5_725 (.A1(n_5_210), .A2(n_5_144), .A3(n_5_713), .ZN(n_5_3975));
   INV_X1 i_5_753 (.A(n_5_444), .ZN(n_5_3976));
   XNOR2_X1 i_5_754 (.A(n_5_4121), .B(m[0]), .ZN(n_5_444));
   XNOR2_X1 i_5_730 (.A(n_5_445), .B(n_5_506), .ZN(n_5_3977));
   NAND2_X1 i_5_745 (.A1(n_5_4113), .A2(n_5_4561), .ZN(n_5_445));
   XOR2_X1 i_5_691 (.A(n_5_4348), .B(n_5_4458), .Z(n_5_3979));
   XNOR2_X1 i_5_534 (.A(n_5_451), .B(n_5_4215), .ZN(n_5_4642));
   NAND2_X1 i_5_541 (.A1(n_5_4207), .A2(n_5_4206), .ZN(n_5_451));
   NAND2_X1 i_5_568 (.A1(n_5_453), .A2(n_5_527), .ZN(n_5_364));
   INV_X1 i_5_738 (.A(n_5_523), .ZN(n_5_453));
   XOR2_X1 i_5_459 (.A(n_5_482), .B(n_5_4321), .Z(n_5_367));
   NAND2_X1 i_5_664 (.A1(n_5_500), .A2(n_5_3996), .ZN(n_5_372));
   NAND2_X1 i_5_769 (.A1(n_5_480), .A2(n_5_4683), .ZN(n_5_373));
   NAND2_X1 i_5_770 (.A1(n_5_481), .A2(n_5_489), .ZN(n_5_480));
   INV_X1 i_5_771 (.A(n_53), .ZN(n_5_4644));
   OAI21_X1 i_5_772 (.A(n_5_490), .B1(n_5_501), .B2(n_5_504), .ZN(n_5_481));
   OAI21_X1 i_5_467 (.A(n_5_4299), .B1(n_5_487), .B2(n_5_4371), .ZN(n_5_482));
   INV_X1 i_5_250 (.A(n_5_4206), .ZN(n_5_483));
   INV_X1 i_5_694 (.A(n_5_4309), .ZN(n_5_3987));
   INV_X1 i_5_520 (.A(n_5_4300), .ZN(n_5_487));
   INV_X1 i_5_777 (.A(n_76), .ZN(n_5_4645));
   INV_X1 i_5_778 (.A(n_61), .ZN(n_5_488));
   NAND2_X1 i_5_779 (.A1(n_5_4361), .A2(n_5_488), .ZN(n_5_489));
   NAND2_X1 i_5_780 (.A1(n_5_4359), .A2(n_61), .ZN(n_5_490));
   NAND2_X1 i_5_781 (.A1(n_5_4361), .A2(n_5_488), .ZN(n_5_3989));
   NAND2_X1 i_5_782 (.A1(n_5_481), .A2(n_5_489), .ZN(n_5_493));
   INV_X1 i_5_783 (.A(n_5_493), .ZN(n_5_495));
   NAND2_X1 i_5_784 (.A1(n_5_4685), .A2(n_5_495), .ZN(n_5_374));
   NAND2_X1 i_5_785 (.A1(n_5_551), .A2(n_5_482), .ZN(n_5_500));
   NAND2_X1 i_5_433 (.A1(n_5_482), .A2(n_5_551), .ZN(n_5_3990));
   AOI22_X1 i_5_787 (.A1(n_5_3990), .A2(n_5_3996), .B1(n_5_548), .B2(n_75), 
      .ZN(n_5_501));
   NOR2_X1 i_5_788 (.A1(n_5_548), .A2(n_75), .ZN(n_5_504));
   INV_X1 i_5_789 (.A(n_75), .ZN(n_5_505));
   NAND2_X1 i_5_452 (.A1(n_5_4407), .A2(n_5_505), .ZN(n_5_3991));
   AOI21_X1 i_5_751 (.A(n_5_4127), .B1(n_5_540), .B2(n_5_541), .ZN(n_5_506));
   INV_X1 i_5_792 (.A(n_5_4127), .ZN(n_5_620));
   NAND2_X1 i_5_793 (.A1(n_5_540), .A2(n_5_541), .ZN(n_5_723));
   OAI21_X1 i_5_253 (.A(n_5_4207), .B1(n_5_4215), .B2(n_5_483), .ZN(n_5_509));
   XOR2_X1 i_5_275 (.A(n_5_4169), .B(n_5_509), .Z(n_5_3993));
   NAND2_X1 i_5_796 (.A1(n_5_513), .A2(n_5_521), .ZN(n_5_510));
   OAI21_X1 i_5_277 (.A(n_5_4207), .B1(n_5_4215), .B2(n_5_483), .ZN(n_5_513));
   NOR2_X1 i_5_798 (.A1(n_5_4762), .A2(n_60), .ZN(n_5_4646));
   INV_X1 i_5_799 (.A(n_60), .ZN(n_5_514));
   NAND2_X1 i_5_800 (.A1(n_5_4762), .A2(n_60), .ZN(n_5_4647));
   INV_X1 i_5_801 (.A(n_60), .ZN(n_5_375));
   INV_X1 i_5_802 (.A(n_5_514), .ZN(n_5_516));
   NAND2_X1 i_5_803 (.A1(n_5_4461), .A2(n_58), .ZN(n_5_3994));
   OR2_X1 i_5_804 (.A1(n_5_4170), .A2(n_69), .ZN(n_5_519));
   NAND2_X1 i_5_805 (.A1(n_5_4170), .A2(n_69), .ZN(n_5_521));
   NOR2_X1 i_5_794 (.A1(n_5_419), .A2(n_55), .ZN(n_5_523));
   NAND2_X1 i_5_807 (.A1(n_5_419), .A2(n_55), .ZN(n_5_527));
   NAND2_X1 i_5_453 (.A1(n_5_4704), .A2(n_5_4645), .ZN(n_5_3996));
   NAND2_X1 i_5_812 (.A1(n_5_510), .A2(n_5_519), .ZN(n_5_4648));
   NAND2_X1 i_5_813 (.A1(n_5_516), .A2(n_5_375), .ZN(n_5_530));
   INV_X1 i_5_814 (.A(n_5_530), .ZN(n_5_376));
   NAND2_X1 i_5_500 (.A1(n_5_537), .A2(n_5_4761), .ZN(n_5_533));
   NAND2_X1 i_5_507 (.A1(n_5_510), .A2(n_5_519), .ZN(n_5_534));
   XNOR2_X1 i_5_526 (.A(n_5_533), .B(n_5_534), .ZN(n_5_377));
   INV_X1 i_5_819 (.A(n_5_4762), .ZN(n_5_535));
   NAND2_X1 i_5_820 (.A1(n_5_535), .A2(n_5_516), .ZN(n_5_537));
   AOI21_X1 i_5_714 (.A(n_5_538), .B1(n_5_3994), .B2(n_5_4348), .ZN(n_5_3998));
   NOR2_X1 i_5_822 (.A1(n_5_4461), .A2(n_58), .ZN(n_5_538));
   NAND2_X1 i_5_823 (.A1(n_5_4159), .A2(n_5_2568), .ZN(n_5_540));
   NAND2_X1 i_5_824 (.A1(n_5_4187), .A2(m[0]), .ZN(n_5_541));
   NAND2_X1 i_5_825 (.A1(n_5_4187), .A2(m[0]), .ZN(n_5_542));
   INV_X1 i_5_826 (.A(n_5_542), .ZN(n_5_543));
   NAND2_X1 i_5_827 (.A1(n_5_4127), .A2(n_5_543), .ZN(n_5_544));
   XNOR2_X1 i_5_828 (.A(n_5_4161), .B(n_5_543), .ZN(n_5_547));
   OAI21_X1 i_5_829 (.A(n_5_544), .B1(n_5_547), .B2(n_5_4127), .ZN(n_5_3999));
   BUF_X1 rt_shieldBuf__2__2__15 (.A(n_5_616), .Z(n_5_548));
   NAND2_X1 i_5_517 (.A1(n_5_4778), .A2(n_76), .ZN(n_5_551));
   NAND2_X1 i_5_831 (.A1(n_5_826), .A2(n_5_420), .ZN(n_5_552));
   NAND2_X1 i_5_832 (.A1(n_5_699), .A2(n_5_378), .ZN(n_5_553));
   NAND2_X1 i_5_833 (.A1(n_5_735), .A2(n_5_4649), .ZN(n_5_555));
   NAND3_X1 i_5_834 (.A1(n_5_552), .A2(n_5_553), .A3(n_5_555), .ZN(n_89));
   NAND2_X1 i_5_482 (.A1(n_5_4278), .A2(n_5_420), .ZN(n_5_4001));
   NAND2_X1 i_5_487 (.A1(n_5_4143), .A2(n_5_378), .ZN(n_5_4002));
   NAND2_X1 i_5_488 (.A1(n_5_293), .A2(n_5_4649), .ZN(n_5_4003));
   INV_X1 i_5_838 (.A(r[6]), .ZN(n_5_560));
   NAND2_X1 i_5_839 (.A1(n_5_718), .A2(n_5_378), .ZN(n_5_566));
   NAND2_X1 i_5_840 (.A1(r[7]), .A2(n_5_560), .ZN(n_5_567));
   NAND2_X1 i_5_841 (.A1(n_5_829), .A2(n_5_420), .ZN(n_5_569));
   XNOR2_X1 i_5_842 (.A(r[7]), .B(r[6]), .ZN(n_5_4649));
   NAND3_X1 i_5_843 (.A1(n_5_566), .A2(n_5_569), .A3(n_5_4015), .ZN(n_5_381));
   NAND2_X1 i_5_844 (.A1(n_5_3795), .A2(n_5_4649), .ZN(n_5_570));
   NAND2_X1 i_5_845 (.A1(n_5_703), .A2(n_5_378), .ZN(n_5_573));
   NAND2_X1 i_5_623 (.A1(n_5_4052), .A2(n_5_4649), .ZN(n_5_724));
   NAND2_X1 i_5_847 (.A1(n_5_3919), .A2(n_5_4649), .ZN(n_5_4005));
   NAND2_X1 i_5_848 (.A1(n_5_4120), .A2(n_5_4649), .ZN(n_5_4006));
   NAND2_X1 i_5_849 (.A1(n_5_870), .A2(n_5_420), .ZN(n_5_4007));
   NAND2_X1 i_5_542 (.A1(n_5_3793), .A2(n_5_4649), .ZN(n_5_574));
   NAND2_X1 i_5_851 (.A1(n_5_917), .A2(n_5_4649), .ZN(n_5_575));
   NAND2_X1 i_5_853 (.A1(n_5_4686), .A2(n_5_4649), .ZN(n_5_410));
   NAND2_X1 i_5_567 (.A1(n_5_850), .A2(n_5_420), .ZN(n_5_418));
   NAND3_X1 i_5_511 (.A1(n_5_4558), .A2(n_5_583), .A3(n_5_582), .ZN(n_5_419));
   NAND2_X1 i_5_608 (.A1(n_5_4188), .A2(n_5_4649), .ZN(n_5_582));
   NAND2_X1 i_5_649 (.A1(n_5_849), .A2(n_5_420), .ZN(n_5_583));
   NAND2_X1 i_5_761 (.A1(n_5_3884), .A2(n_5_4649), .ZN(n_5_4010));
   NAND2_X1 i_5_768 (.A1(n_5_838), .A2(n_5_420), .ZN(n_5_4011));
   NAND2_X1 i_5_857 (.A1(n_5_930), .A2(n_5_378), .ZN(n_5_4012));
   NAND2_X1 i_5_861 (.A1(n_5_828), .A2(n_5_420), .ZN(n_5_4013));
   INV_X1 i_5_862 (.A(n_5_567), .ZN(n_5_420));
   NOR2_X1 i_5_863 (.A1(r[7]), .A2(n_5_560), .ZN(n_5_378));
   NAND2_X1 i_5_864 (.A1(n_5_3727), .A2(n_5_4649), .ZN(n_5_4015));
   NAND2_X1 i_5_865 (.A1(n_5_3672), .A2(n_5_4017), .ZN(n_5_584));
   NAND2_X1 i_5_866 (.A1(n_5_3142), .A2(n_5_3333), .ZN(n_5_585));
   NAND2_X1 i_5_867 (.A1(n_5_3365), .A2(n_5_599), .ZN(n_5_586));
   NAND3_X1 i_5_868 (.A1(n_5_584), .A2(n_5_585), .A3(n_5_586), .ZN(n_5_587));
   NAND2_X1 i_5_869 (.A1(n_5_3381), .A2(n_5_599), .ZN(n_5_588));
   NAND2_X1 i_5_870 (.A1(n_5_3401), .A2(n_5_599), .ZN(n_5_589));
   NAND2_X1 i_5_871 (.A1(n_5_4192), .A2(n_5_599), .ZN(n_5_593));
   INV_X1 i_5_872 (.A(n_5_593), .ZN(n_5_3332));
   NAND2_X1 i_5_873 (.A1(n_5_4108), .A2(n_5_599), .ZN(n_5_595));
   INV_X1 i_5_874 (.A(r[5]), .ZN(n_5_596));
   NAND2_X1 i_5_875 (.A1(r[6]), .A2(n_5_596), .ZN(n_5_598));
   XNOR2_X1 i_5_876 (.A(r[6]), .B(r[5]), .ZN(n_5_599));
   INV_X1 i_5_877 (.A(n_5_600), .ZN(n_5_3333));
   NAND2_X1 i_5_878 (.A1(n_5_601), .A2(n_5_604), .ZN(n_5_600));
   NAND2_X1 i_5_879 (.A1(n_5_3372), .A2(n_5_599), .ZN(n_5_4653));
   INV_X1 i_5_880 (.A(r[6]), .ZN(n_5_601));
   INV_X1 i_5_881 (.A(n_5_596), .ZN(n_5_604));
   NAND2_X1 i_5_882 (.A1(n_5_599), .A2(n_5_4101), .ZN(n_5_605));
   NAND2_X1 i_5_883 (.A1(n_5_3578), .A2(n_5_4017), .ZN(n_5_606));
   NAND2_X1 i_5_884 (.A1(n_5_3152), .A2(n_5_1006), .ZN(n_5_611));
   INV_X1 i_5_885 (.A(r[6]), .ZN(n_5_612));
   NAND2_X1 i_5_886 (.A1(n_5_4140), .A2(n_5_599), .ZN(n_5_4016));
   NAND2_X1 i_5_575 (.A1(n_5_4155), .A2(n_5_599), .ZN(n_5_613));
   NAND3_X1 i_5_512 (.A1(n_5_615), .A2(n_5_618), .A3(n_5_614), .ZN(n_5_293));
   NAND2_X1 i_5_603 (.A1(n_5_678), .A2(n_5_599), .ZN(n_5_614));
   NAND2_X1 i_5_513 (.A1(n_5_3878), .A2(n_5_4017), .ZN(n_5_615));
   NAND2_X1 i_5_522 (.A1(n_5_3147), .A2(n_5_1006), .ZN(n_5_618));
   NAND2_X1 i_5_892 (.A1(n_5_3377), .A2(n_5_599), .ZN(n_5_621));
   NAND2_X1 i_5_893 (.A1(n_5_4512), .A2(n_5_4017), .ZN(n_5_436));
   NAND2_X1 i_5_894 (.A1(n_5_3148), .A2(n_5_1006), .ZN(n_5_623));
   INV_X1 i_5_895 (.A(n_5_598), .ZN(n_5_4017));
   NAND2_X1 i_5_896 (.A1(n_5_3399), .A2(n_5_599), .ZN(n_5_3335));
   NOR2_X1 i_5_897 (.A1(r[6]), .A2(n_5_596), .ZN(n_5_1006));
   NAND2_X1 i_5_898 (.A1(n_5_612), .A2(r[5]), .ZN(n_5_624));
   INV_X1 i_5_899 (.A(n_5_624), .ZN(n_5_635));
   NAND2_X1 i_5_900 (.A1(n_5_601), .A2(n_5_604), .ZN(n_5_637));
   INV_X1 i_5_901 (.A(n_5_637), .ZN(n_5_638));
   NAND2_X1 i_5_902 (.A1(n_5_612), .A2(r[5]), .ZN(n_5_639));
   INV_X1 i_5_903 (.A(n_5_639), .ZN(n_5_640));
   NAND2_X1 i_5_904 (.A1(n_5_4150), .A2(n_5_599), .ZN(n_5_4019));
   NAND2_X1 i_5_905 (.A1(n_5_612), .A2(r[5]), .ZN(n_5_641));
   INV_X1 i_5_906 (.A(n_5_641), .ZN(n_5_3338));
   NAND2_X1 i_5_907 (.A1(n_5_3983), .A2(n_5_599), .ZN(n_5_4020));
   NAND2_X1 i_5_659 (.A1(n_5_3829), .A2(n_5_4017), .ZN(n_5_643));
   INV_X1 i_5_665 (.A(n_5_589), .ZN(n_5_644));
   AOI21_X1 i_5_667 (.A(n_5_644), .B1(n_5_3151), .B2(n_5_638), .ZN(n_5_645));
   INV_X1 i_5_911 (.A(n_5_588), .ZN(n_5_648));
   AOI21_X1 i_5_912 (.A(n_5_648), .B1(n_5_3581), .B2(n_5_4017), .ZN(n_5_652));
   INV_X1 i_5_591 (.A(n_5_613), .ZN(n_5_653));
   NAND2_X1 i_5_914 (.A1(n_5_612), .A2(r[5]), .ZN(n_5_654));
   INV_X1 i_5_915 (.A(n_5_654), .ZN(n_5_665));
   NAND2_X1 i_5_916 (.A1(n_5_3160), .A2(n_5_665), .ZN(n_5_667));
   INV_X1 i_5_917 (.A(m[14]), .ZN(n_5_669));
   INV_X1 i_5_918 (.A(m[15]), .ZN(n_5_672));
   NAND2_X1 i_5_919 (.A1(n_5_587), .A2(m[0]), .ZN(n_5_673));
   INV_X1 i_5_920 (.A(m[1]), .ZN(n_5_4021));
   INV_X1 i_5_921 (.A(m[2]), .ZN(n_5_674));
   INV_X1 i_5_922 (.A(m[13]), .ZN(n_5_676));
   NAND2_X1 i_5_923 (.A1(n_5_3727), .A2(m[14]), .ZN(n_5_677));
   INV_X1 i_5_924 (.A(n_5_3727), .ZN(n_5_680));
   NAND2_X1 i_5_925 (.A1(n_5_825), .A2(n_5_815), .ZN(n_5_681));
   OAI21_X1 i_5_926 (.A(n_5_815), .B1(n_5_4275), .B2(n_5_673), .ZN(n_5_3124));
   NAND2_X1 i_5_927 (.A1(n_5_915), .A2(n_5_4270), .ZN(n_5_689));
   NAND2_X1 i_5_547 (.A1(n_5_704), .A2(n_5_4414), .ZN(n_5_4022));
   NAND3_X1 i_5_929 (.A1(n_5_752), .A2(n_5_4025), .A3(n_5_755), .ZN(n_5_691));
   NAND2_X1 i_5_930 (.A1(n_5_677), .A2(n_5_738), .ZN(n_5_695));
   NAND2_X1 i_5_931 (.A1(n_5_695), .A2(n_5_4025), .ZN(n_5_697));
   INV_X1 i_5_932 (.A(m[0]), .ZN(n_5_698));
   XNOR2_X1 i_5_933 (.A(n_5_735), .B(n_5_698), .ZN(n_5_699));
   XNOR2_X1 i_5_934 (.A(n_5_3798), .B(n_5_814), .ZN(n_5_703));
   XNOR2_X1 i_5_936 (.A(n_5_3727), .B(m[14]), .ZN(n_5_3339));
   INV_X1 i_5_565 (.A(n_5_4270), .ZN(n_5_704));
   OAI211_X1 i_5_938 (.A(n_5_743), .B(n_5_3770), .C1(n_5_707), .C2(n_5_706), 
      .ZN(n_5_705));
   NAND2_X1 i_5_939 (.A1(n_5_798), .A2(n_5_4238), .ZN(n_5_706));
   AND2_X1 i_5_940 (.A1(n_5_794), .A2(n_5_3762), .ZN(n_5_707));
   OAI21_X1 i_5_592 (.A(n_5_915), .B1(n_5_797), .B2(n_5_4269), .ZN(n_5_708));
   NAND3_X1 i_5_544 (.A1(n_5_714), .A2(n_5_440), .A3(n_5_4415), .ZN(n_5_709));
   OAI21_X1 i_5_548 (.A(n_5_4270), .B1(n_5_4023), .B2(n_5_715), .ZN(n_5_714));
   INV_X1 i_5_555 (.A(n_5_4414), .ZN(n_5_715));
   AND2_X1 i_5_577 (.A1(n_5_797), .A2(n_5_915), .ZN(n_5_4023));
   INV_X1 i_5_946 (.A(m[9]), .ZN(n_5_4024));
   XNOR2_X1 i_5_566 (.A(n_5_4719), .B(n_5_3515), .ZN(n_5_438));
   NAND3_X1 i_5_948 (.A1(n_5_4548), .A2(n_5_754), .A3(n_5_4549), .ZN(n_5_717));
   NAND2_X1 i_5_949 (.A1(n_5_720), .A2(n_5_719), .ZN(n_5_718));
   NAND3_X1 i_5_950 (.A1(n_5_750), .A2(n_5_726), .A3(n_5_722), .ZN(n_5_719));
   NAND2_X1 i_5_951 (.A1(n_5_725), .A2(n_5_721), .ZN(n_5_720));
   INV_X1 i_5_952 (.A(n_5_722), .ZN(n_5_721));
   XNOR2_X1 i_5_953 (.A(m[14]), .B(n_5_672), .ZN(n_5_722));
   NAND2_X1 i_5_954 (.A1(n_5_750), .A2(n_5_726), .ZN(n_5_725));
   INV_X1 i_5_955 (.A(n_5_727), .ZN(n_5_726));
   NAND2_X1 i_5_956 (.A1(n_5_691), .A2(n_5_697), .ZN(n_5_727));
   OAI21_X1 i_5_586 (.A(n_5_911), .B1(n_5_729), .B2(n_5_4454), .ZN(n_5_439));
   AOI21_X1 i_5_604 (.A(n_5_689), .B1(n_5_791), .B2(n_5_792), .ZN(n_5_729));
   AOI21_X1 i_5_960 (.A(n_5_818), .B1(n_5_3761), .B2(n_5_3762), .ZN(n_5_3126));
   INV_X1 i_5_961 (.A(m[4]), .ZN(n_5_730));
   INV_X1 i_5_962 (.A(n_5_4052), .ZN(n_5_731));
   INV_X1 i_5_963 (.A(m[3]), .ZN(n_5_732));
   INV_X1 i_5_964 (.A(m[5]), .ZN(n_5_3340));
   INV_X1 i_5_965 (.A(m[7]), .ZN(n_5_733));
   NAND2_X1 i_5_966 (.A1(n_5_669), .A2(n_5_680), .ZN(n_5_4025));
   INV_X1 i_5_967 (.A(m[12]), .ZN(n_5_734));
   BUF_X1 rt_shieldBuf__2__2__3 (.A(n_5_587), .Z(n_5_735));
   INV_X1 i_5_968 (.A(m[1]), .ZN(n_5_736));
   XNOR2_X1 i_5_969 (.A(n_5_3562), .B(n_5_673), .ZN(n_5_737));
   INV_X1 i_5_970 (.A(n_5_734), .ZN(n_5_3128));
   NAND2_X1 i_5_971 (.A1(n_5_753), .A2(n_5_676), .ZN(n_5_738));
   NAND2_X1 i_5_644 (.A1(m[10]), .A2(n_5_4188), .ZN(n_5_440));
   INV_X1 i_5_973 (.A(n_5_793), .ZN(n_5_3129));
   INV_X1 i_5_974 (.A(n_5_733), .ZN(n_5_740));
   NAND2_X1 i_5_975 (.A1(n_5_4053), .A2(n_5_4024), .ZN(n_5_741));
   NAND2_X1 i_5_976 (.A1(n_5_741), .A2(n_5_4688), .ZN(n_5_742));
   NAND2_X1 i_5_977 (.A1(m[5]), .A2(n_5_4120), .ZN(n_5_743));
   NAND2_X1 i_5_978 (.A1(n_5_755), .A2(n_5_754), .ZN(n_5_744));
   INV_X1 i_5_979 (.A(n_5_744), .ZN(n_5_4026));
   NAND2_X1 i_5_980 (.A1(n_5_4029), .A2(n_5_717), .ZN(n_5_745));
   NAND2_X1 i_5_981 (.A1(n_5_4167), .A2(n_5_3340), .ZN(n_5_4027));
   NAND2_X1 i_5_982 (.A1(n_5_4167), .A2(n_5_3340), .ZN(n_5_4028));
   XNOR2_X1 i_5_653 (.A(n_5_293), .B(m[11]), .ZN(n_5_746));
   NAND2_X1 i_5_984 (.A1(n_5_4548), .A2(n_5_4549), .ZN(n_5_747));
   INV_X1 i_5_985 (.A(n_5_747), .ZN(n_5_748));
   NAND2_X1 i_5_986 (.A1(n_5_4389), .A2(n_5_748), .ZN(n_5_750));
   INV_X1 i_5_987 (.A(m[13]), .ZN(n_5_751));
   INV_X1 i_5_988 (.A(n_5_4029), .ZN(n_5_752));
   INV_X1 i_5_989 (.A(n_5_3884), .ZN(n_5_753));
   NAND2_X1 i_5_990 (.A1(n_5_734), .A2(n_5_4787), .ZN(n_5_4029));
   NAND2_X1 i_5_991 (.A1(m[12]), .A2(n_5_3933), .ZN(n_5_754));
   NAND2_X1 i_5_992 (.A1(m[13]), .A2(n_5_3884), .ZN(n_5_755));
   NAND2_X1 i_5_993 (.A1(n_5_4668), .A2(n_5_4691), .ZN(n_5_756));
   NAND2_X1 i_5_994 (.A1(n_5_3933), .A2(m[12]), .ZN(n_5_757));
   INV_X1 i_5_995 (.A(m[13]), .ZN(n_5_758));
   NAND2_X1 i_5_996 (.A1(n_5_4549), .A2(n_5_758), .ZN(n_5_759));
   INV_X1 i_5_997 (.A(n_5_759), .ZN(n_5_760));
   NAND2_X1 i_5_998 (.A1(n_5_734), .A2(n_5_758), .ZN(n_5_761));
   INV_X1 i_5_999 (.A(n_5_761), .ZN(n_5_762));
   INV_X1 i_5_1000 (.A(n_5_676), .ZN(n_5_763));
   NAND3_X1 i_5_1001 (.A1(n_5_4668), .A2(n_5_4691), .A3(n_5_763), .ZN(n_5_764));
   INV_X1 i_5_1002 (.A(m[12]), .ZN(n_5_765));
   NOR2_X1 i_5_1003 (.A1(n_5_676), .A2(n_5_765), .ZN(n_5_766));
   NAND2_X1 i_5_1004 (.A1(n_5_3933), .A2(n_5_766), .ZN(n_5_767));
   INV_X1 i_5_1005 (.A(n_5_4549), .ZN(n_5_768));
   NAND2_X1 i_5_1006 (.A1(n_5_768), .A2(n_5_763), .ZN(n_5_769));
   NAND3_X1 i_5_1007 (.A1(n_5_764), .A2(n_5_767), .A3(n_5_769), .ZN(n_5_770));
   NAND2_X1 i_5_1008 (.A1(n_5_4787), .A2(n_5_734), .ZN(n_5_771));
   NAND2_X1 i_5_1009 (.A1(n_5_770), .A2(n_5_771), .ZN(n_5_772));
   NAND2_X1 i_5_1010 (.A1(n_5_3894), .A2(n_5_772), .ZN(n_5_3341));
   INV_X1 i_5_1011 (.A(n_5_681), .ZN(n_5_773));
   AOI21_X1 i_5_673 (.A(n_5_3778), .B1(n_5_3507), .B2(n_5_773), .ZN(n_5_4030));
   NAND2_X1 i_5_1013 (.A1(n_5_4414), .A2(n_5_788), .ZN(n_5_4031));
   NAND2_X1 i_5_1014 (.A1(n_5_733), .A2(n_5_4498), .ZN(n_5_774));
   INV_X1 i_5_1015 (.A(m[7]), .ZN(n_5_775));
   INV_X1 i_5_1016 (.A(n_5_733), .ZN(n_5_776));
   INV_X1 i_5_1017 (.A(m[6]), .ZN(n_5_777));
   NAND2_X1 i_5_1018 (.A1(n_5_777), .A2(n_5_733), .ZN(n_5_778));
   INV_X1 i_5_1019 (.A(n_5_733), .ZN(n_5_779));
   NAND2_X1 i_5_1020 (.A1(n_5_778), .A2(n_5_779), .ZN(n_5_780));
   INV_X1 i_5_1021 (.A(n_5_780), .ZN(n_5_781));
   AOI21_X1 i_5_1022 (.A(n_5_781), .B1(n_5_4694), .B2(n_5_778), .ZN(n_5_782));
   NAND2_X1 i_5_1023 (.A1(n_5_933), .A2(n_5_782), .ZN(n_5_783));
   INV_X1 i_5_1024 (.A(n_5_933), .ZN(n_5_784));
   INV_X1 i_5_1026 (.A(m[11]), .ZN(n_5_785));
   XNOR2_X1 i_5_668 (.A(n_5_293), .B(n_5_785), .ZN(n_5_786));
   NAND2_X1 i_5_669 (.A1(n_5_709), .A2(n_5_911), .ZN(n_5_787));
   NAND2_X1 i_5_1029 (.A1(m[8]), .A2(n_5_917), .ZN(n_5_788));
   NAND2_X1 i_5_1030 (.A1(n_5_917), .A2(m[8]), .ZN(n_5_4032));
   NAND2_X1 i_5_1031 (.A1(n_5_4018), .A2(n_5_730), .ZN(n_5_789));
   NAND2_X1 i_5_1032 (.A1(n_5_3919), .A2(m[4]), .ZN(n_5_790));
   NAND2_X1 i_5_1033 (.A1(n_5_789), .A2(n_5_790), .ZN(n_5_3131));
   NAND2_X1 i_5_1034 (.A1(n_5_774), .A2(n_5_3538), .ZN(n_5_791));
   OAI21_X1 i_5_1035 (.A(n_5_783), .B1(n_5_3793), .B2(n_5_784), .ZN(n_5_792));
   NAND2_X1 i_5_1036 (.A1(n_5_4120), .A2(m[5]), .ZN(n_5_793));
   INV_X1 i_5_1037 (.A(n_5_4118), .ZN(n_5_4033));
   NAND2_X1 i_5_1038 (.A1(n_5_3343), .A2(n_5_4175), .ZN(n_5_794));
   NAND2_X1 i_5_1039 (.A1(n_5_3538), .A2(n_5_774), .ZN(n_5_795));
   OAI21_X1 i_5_1040 (.A(n_5_783), .B1(n_5_784), .B2(n_5_3793), .ZN(n_5_796));
   NAND2_X1 i_5_1041 (.A1(n_5_795), .A2(n_5_796), .ZN(n_5_797));
   NAND2_X1 i_5_1042 (.A1(n_5_3340), .A2(n_5_4167), .ZN(n_5_798));
   NAND3_X1 i_5_1043 (.A1(n_5_4014), .A2(n_5_4004), .A3(n_5_4016), .ZN(n_5_799));
   INV_X1 i_5_1044 (.A(n_5_799), .ZN(n_5_800));
   INV_X1 i_5_1045 (.A(n_5_776), .ZN(n_5_801));
   NAND2_X1 i_5_1046 (.A1(n_5_800), .A2(n_5_801), .ZN(n_5_802));
   INV_X1 i_5_1047 (.A(n_5_775), .ZN(n_5_803));
   NAND2_X1 i_5_1048 (.A1(n_5_799), .A2(n_5_803), .ZN(n_5_804));
   NAND2_X1 i_5_1049 (.A1(n_5_705), .A2(n_5_3494), .ZN(n_5_805));
   INV_X1 i_5_1050 (.A(n_5_378), .ZN(n_5_806));
   NAND4_X1 i_5_569 (.A1(n_5_805), .A2(n_5_802), .A3(n_5_804), .A4(n_5_378), 
      .ZN(n_5_807));
   NAND2_X1 i_5_572 (.A1(n_5_4191), .A2(n_5_807), .ZN(n_5_808));
   INV_X1 i_5_580 (.A(n_5_574), .ZN(n_5_809));
   NOR2_X1 i_5_595 (.A1(n_5_808), .A2(n_5_809), .ZN(n_5_4034));
   NAND2_X1 i_5_1055 (.A1(n_5_4273), .A2(n_5_4021), .ZN(n_5_810));
   NAND2_X1 i_5_1056 (.A1(n_5_816), .A2(n_5_810), .ZN(n_5_811));
   INV_X1 i_5_1057 (.A(n_5_673), .ZN(n_5_812));
   NAND2_X1 i_5_1058 (.A1(n_5_810), .A2(n_5_812), .ZN(n_5_813));
   NAND2_X1 i_5_1059 (.A1(n_5_811), .A2(n_5_813), .ZN(n_5_814));
   NAND3_X1 i_5_1060 (.A1(n_5_3506), .A2(n_5_3507), .A3(n_5_3505), .ZN(n_5_3343));
   NAND2_X1 i_5_1061 (.A1(n_5_3563), .A2(m[1]), .ZN(n_5_815));
   INV_X1 i_5_1062 (.A(n_5_3561), .ZN(n_5_816));
   INV_X1 i_5_1063 (.A(n_5_3340), .ZN(n_5_817));
   NOR2_X1 i_5_1064 (.A1(n_5_4120), .A2(n_5_817), .ZN(n_5_818));
   INV_X1 i_5_658 (.A(n_5_742), .ZN(n_5_819));
   XNOR2_X1 i_5_678 (.A(n_5_819), .B(n_5_708), .ZN(n_5_820));
   NAND2_X1 i_5_680 (.A1(n_5_820), .A2(n_5_378), .ZN(n_5_452));
   NAND2_X1 i_5_1068 (.A1(n_5_601), .A2(n_5_604), .ZN(n_5_822));
   INV_X1 i_5_1069 (.A(n_5_822), .ZN(n_5_3345));
   NAND2_X1 i_5_1070 (.A1(n_5_4273), .A2(n_5_4021), .ZN(n_5_823));
   INV_X1 i_5_1071 (.A(n_5_673), .ZN(n_5_824));
   NAND2_X1 i_5_1072 (.A1(n_5_823), .A2(n_5_824), .ZN(n_5_825));
   INV_X1 i_5_1073 (.A(n_5_827), .ZN(n_5_826));
   OAI21_X1 i_5_1074 (.A(n_5_891), .B1(m[0]), .B2(n_5_735), .ZN(n_5_827));
   XNOR2_X1 i_5_1075 (.A(n_5_886), .B(n_5_922), .ZN(n_5_828));
   XNOR2_X1 i_5_1076 (.A(n_5_831), .B(n_5_830), .ZN(n_5_829));
   XNOR2_X1 i_5_1077 (.A(n_54), .B(n_53), .ZN(n_5_830));
   AOI21_X1 i_5_1078 (.A(n_5_865), .B1(n_5_833), .B2(n_5_832), .ZN(n_5_831));
   INV_X1 i_5_1079 (.A(n_5_3727), .ZN(n_5_832));
   INV_X1 i_5_1080 (.A(n_53), .ZN(n_5_833));
   INV_X1 i_5_1081 (.A(n_75), .ZN(n_5_834));
   INV_X1 i_5_810 (.A(n_5_293), .ZN(n_5_835));
   INV_X1 i_5_1083 (.A(n_76), .ZN(n_5_836));
   NAND2_X1 i_5_597 (.A1(n_5_3735), .A2(n_5_3769), .ZN(n_5_837));
   NAND2_X1 i_5_835 (.A1(n_5_835), .A2(n_5_836), .ZN(n_5_4035));
   NAND2_X1 i_5_858 (.A1(n_5_3840), .A2(n_5_890), .ZN(n_5_838));
   INV_X1 i_5_1087 (.A(n_5_3933), .ZN(n_5_839));
   INV_X1 i_5_1088 (.A(n_75), .ZN(n_5_840));
   INV_X1 i_5_1089 (.A(n_5_3185), .ZN(n_5_841));
   INV_X1 i_5_1090 (.A(n_73), .ZN(n_5_4036));
   INV_X1 i_5_1091 (.A(n_61), .ZN(n_5_387));
   OAI21_X1 i_5_672 (.A(n_5_856), .B1(n_5_851), .B2(n_5_857), .ZN(n_5_844));
   NAND2_X1 i_5_889 (.A1(n_5_4366), .A2(n_5_844), .ZN(n_5_845));
   NAND3_X1 i_5_1096 (.A1(n_5_845), .A2(n_5_4790), .A3(n_5_912), .ZN(n_5_846));
   OAI21_X1 i_5_609 (.A(n_5_837), .B1(n_5_3185), .B2(n_5_4694), .ZN(n_5_847));
   NAND2_X1 i_5_683 (.A1(n_5_4366), .A2(n_5_912), .ZN(n_5_848));
   XNOR2_X1 i_5_762 (.A(n_5_848), .B(n_5_844), .ZN(n_5_849));
   NAND2_X1 i_5_677 (.A1(n_5_845), .A2(n_5_912), .ZN(n_5_4038));
   INV_X1 i_5_891 (.A(n_5_4038), .ZN(n_5_4039));
   XOR2_X1 i_5_684 (.A(n_5_899), .B(n_5_908), .Z(n_5_850));
   AOI21_X1 i_5_1103 (.A(n_5_869), .B1(n_5_900), .B2(n_5_3986), .ZN(n_5_851));
   NAND2_X1 i_5_1105 (.A1(n_5_4694), .A2(n_5_3185), .ZN(n_5_852));
   INV_X1 i_5_1106 (.A(n_5_852), .ZN(n_5_853));
   NOR2_X1 i_5_739 (.A1(n_5_904), .A2(n_5_853), .ZN(n_5_854));
   NAND2_X1 i_5_1108 (.A1(n_5_3797), .A2(n_5_906), .ZN(n_5_3136));
   INV_X1 i_5_1109 (.A(n_60), .ZN(n_5_855));
   NAND2_X1 i_5_1110 (.A1(n_5_4686), .A2(n_55), .ZN(n_5_856));
   NOR2_X1 i_5_1111 (.A1(n_5_4686), .A2(n_55), .ZN(n_5_857));
   XNOR2_X1 i_5_1112 (.A(n_5_3919), .B(n_58), .ZN(n_5_3347));
   NAND2_X1 i_5_617 (.A1(n_5_4400), .A2(n_5_4233), .ZN(n_5_858));
   NAND2_X1 i_5_1114 (.A1(n_5_839), .A2(n_5_840), .ZN(n_5_4041));
   NAND2_X1 i_5_746 (.A1(n_5_3793), .A2(n_69), .ZN(n_5_859));
   OAI21_X1 i_5_1116 (.A(n_5_862), .B1(n_5_887), .B2(n_5_877), .ZN(n_5_860));
   XNOR2_X1 i_5_1117 (.A(n_5_4282), .B(n_5_3768), .ZN(n_5_4655));
   INV_X1 i_5_622 (.A(n_5_4232), .ZN(n_5_4042));
   INV_X1 i_5_1119 (.A(n_5_2568), .ZN(n_5_861));
   NAND2_X1 i_5_1120 (.A1(n_5_871), .A2(n_5_879), .ZN(n_5_862));
   NAND2_X1 i_5_1121 (.A1(n_5_3727), .A2(n_53), .ZN(n_5_863));
   NAND2_X1 i_5_1122 (.A1(n_5_924), .A2(n_5_863), .ZN(n_5_864));
   NOR2_X1 i_5_1123 (.A1(n_5_860), .A2(n_5_864), .ZN(n_5_865));
   AOI21_X1 i_5_1124 (.A(n_5_3797), .B1(n_5_902), .B2(n_5_3796), .ZN(n_5_4043));
   AOI21_X1 i_5_696 (.A(n_5_3797), .B1(n_5_902), .B2(n_5_3796), .ZN(n_5_866));
   NAND2_X1 i_5_1126 (.A1(n_5_3557), .A2(n_5_861), .ZN(n_5_867));
   INV_X1 i_5_1127 (.A(n_58), .ZN(n_5_868));
   NAND2_X1 i_5_628 (.A1(n_5_3926), .A2(n_5_868), .ZN(n_5_4044));
   INV_X1 i_5_765 (.A(n_5_914), .ZN(n_5_869));
   XNOR2_X1 i_5_1130 (.A(n_5_3782), .B(n_5_910), .ZN(n_5_870));
   INV_X1 i_5_1131 (.A(n_5_888), .ZN(n_5_871));
   NAND2_X1 i_5_1132 (.A1(n_5_839), .A2(n_5_840), .ZN(n_5_872));
   NAND2_X1 i_5_1133 (.A1(n_5_3981), .A2(n_5_834), .ZN(n_5_3682));
   NAND3_X1 i_5_1134 (.A1(n_5_3808), .A2(n_5_3786), .A3(n_5_3736), .ZN(n_5_421));
   NAND2_X1 i_5_1135 (.A1(n_5_3981), .A2(n_5_834), .ZN(n_5_874));
   INV_X1 i_5_1136 (.A(n_5_874), .ZN(n_5_875));
   NAND2_X1 i_5_1137 (.A1(n_5_875), .A2(n_5_3786), .ZN(n_5_602));
   NOR2_X1 i_5_663 (.A1(n_5_866), .A2(n_5_858), .ZN(n_5_4045));
   INV_X1 i_5_1139 (.A(n_5_879), .ZN(n_5_877));
   INV_X1 i_5_1140 (.A(n_5_3884), .ZN(n_5_842));
   NAND2_X1 i_5_1141 (.A1(n_5_3884), .A2(n_61), .ZN(n_5_879));
   NAND2_X1 i_5_1142 (.A1(n_5_3933), .A2(n_75), .ZN(n_5_3736));
   NAND2_X1 i_5_1143 (.A1(n_5_846), .A2(n_5_4579), .ZN(n_5_3808));
   NAND2_X1 i_5_1144 (.A1(n_5_3787), .A2(n_5_387), .ZN(n_5_880));
   NAND2_X1 i_5_1145 (.A1(n_5_3933), .A2(n_75), .ZN(n_5_881));
   NAND2_X1 i_5_1146 (.A1(n_5_846), .A2(n_5_4579), .ZN(n_5_882));
   NAND2_X1 i_5_1147 (.A1(n_5_881), .A2(n_5_882), .ZN(n_5_883));
   NAND3_X1 i_5_1148 (.A1(n_5_880), .A2(n_5_872), .A3(n_5_883), .ZN(n_5_884));
   NAND2_X1 i_5_1149 (.A1(n_5_3884), .A2(n_61), .ZN(n_5_885));
   NAND2_X1 i_5_1150 (.A1(n_5_884), .A2(n_5_885), .ZN(n_5_886));
   NAND2_X1 i_5_1151 (.A1(n_5_3736), .A2(n_5_3808), .ZN(n_5_887));
   NAND2_X1 i_5_1152 (.A1(n_5_839), .A2(n_5_840), .ZN(n_5_888));
   AOI22_X1 i_5_1153 (.A1(n_5_3808), .A2(n_5_3736), .B1(n_5_839), .B2(n_5_840), 
      .ZN(n_5_889));
   NAND2_X1 i_5_859 (.A1(n_5_921), .A2(n_5_889), .ZN(n_5_890));
   NAND2_X1 i_5_1155 (.A1(n_5_587), .A2(m[0]), .ZN(n_5_891));
   INV_X1 i_5_1156 (.A(n_5_867), .ZN(n_5_892));
   NAND2_X1 i_5_1157 (.A1(n_5_587), .A2(m[0]), .ZN(n_5_893));
   INV_X1 i_5_1158 (.A(n_5_893), .ZN(n_5_894));
   NAND2_X1 i_5_1159 (.A1(n_5_892), .A2(n_5_894), .ZN(n_5_895));
   XNOR2_X1 i_5_1160 (.A(n_5_3558), .B(n_5_894), .ZN(n_5_896));
   OAI21_X1 i_5_1161 (.A(n_5_895), .B1(n_5_896), .B2(n_5_892), .ZN(n_5_897));
   OAI21_X1 i_5_766 (.A(n_5_859), .B1(n_5_854), .B2(n_5_3792), .ZN(n_5_898));
   AOI21_X1 i_5_774 (.A(n_5_869), .B1(n_5_898), .B2(n_5_3986), .ZN(n_5_899));
   OAI21_X1 i_5_1164 (.A(n_5_859), .B1(n_5_854), .B2(n_5_3792), .ZN(n_5_900));
   NAND2_X1 i_5_720 (.A1(n_5_3560), .A2(n_5_891), .ZN(n_5_901));
   NAND2_X1 i_5_734 (.A1(n_5_901), .A2(n_5_927), .ZN(n_5_902));
   NOR2_X1 i_5_1167 (.A1(n_5_4323), .A2(n_5_3352), .ZN(n_5_903));
   NAND2_X1 i_5_1168 (.A1(n_5_4696), .A2(n_5_841), .ZN(n_5_3350));
   NOR2_X1 i_5_1169 (.A1(n_5_903), .A2(n_5_3734), .ZN(n_5_904));
   INV_X1 i_5_1170 (.A(n_69), .ZN(n_5_4048));
   INV_X1 i_5_1171 (.A(n_5_4120), .ZN(n_5_4049));
   INV_X1 i_5_1172 (.A(n_66), .ZN(n_5_4050));
   AOI21_X1 i_5_1173 (.A(n_5_3559), .B1(n_5_3560), .B2(n_5_891), .ZN(n_5_905));
   XNOR2_X1 i_5_1174 (.A(n_5_3796), .B(n_5_905), .ZN(n_5_3138));
   AOI21_X1 i_5_1175 (.A(n_5_3559), .B1(n_5_3560), .B2(n_5_891), .ZN(n_5_906));
   NAND2_X1 i_5_744 (.A1(n_5_643), .A2(n_5_645), .ZN(n_5_3139));
   XNOR2_X1 i_5_752 (.A(n_5_3139), .B(m[3]), .ZN(n_5_4051));
   XNOR2_X1 i_5_755 (.A(n_5_3139), .B(n_65), .ZN(n_5_907));
   NAND2_X1 i_5_756 (.A1(n_5_643), .A2(n_5_645), .ZN(n_5_4052));
   INV_X1 i_5_748 (.A(n_5_3569), .ZN(n_5_4053));
   XNOR2_X1 i_5_776 (.A(n_5_3569), .B(n_55), .ZN(n_5_908));
   NAND3_X1 i_5_679 (.A1(n_5_4202), .A2(n_5_4393), .A3(n_5_3719), .ZN(n_5_909));
   XNOR2_X1 i_5_1183 (.A(n_5_909), .B(n_66), .ZN(n_5_910));
   XNOR2_X1 i_5_688 (.A(n_5_909), .B(n_66), .ZN(n_5_3352));
   OR2_X1 i_5_671 (.A1(m[10]), .A2(n_5_4428), .ZN(n_5_911));
   XNOR2_X1 i_5_763 (.A(n_5_4428), .B(m[10]), .ZN(n_5_455));
   NAND2_X1 i_5_1085 (.A1(n_5_4428), .A2(n_73), .ZN(n_5_912));
   NAND3_X1 i_5_1188 (.A1(n_5_667), .A2(n_5_3729), .A3(n_5_595), .ZN(n_5_913));
   NAND2_X1 i_5_786 (.A1(n_5_917), .A2(n_60), .ZN(n_5_914));
   OR2_X1 i_5_1190 (.A1(m[8]), .A2(n_5_917), .ZN(n_5_915));
   XNOR2_X1 i_5_1191 (.A(n_5_913), .B(m[8]), .ZN(n_5_916));
   NAND3_X1 i_5_1192 (.A1(n_5_667), .A2(n_5_3729), .A3(n_5_595), .ZN(n_5_917));
   NAND2_X1 i_5_1193 (.A1(n_5_3884), .A2(n_61), .ZN(n_5_918));
   INV_X1 i_5_1194 (.A(n_5_842), .ZN(n_5_919));
   INV_X1 i_5_1195 (.A(n_5_387), .ZN(n_5_920));
   OAI21_X1 i_5_1196 (.A(n_5_918), .B1(n_5_919), .B2(n_5_920), .ZN(n_5_921));
   OAI22_X1 i_5_1197 (.A1(n_5_832), .A2(n_5_833), .B1(n_5_3727), .B2(n_53), 
      .ZN(n_5_922));
   NAND2_X1 i_5_1198 (.A1(n_5_4158), .A2(n_5_378), .ZN(n_5_4056));
   NAND2_X1 i_5_1199 (.A1(n_5_731), .A2(n_5_732), .ZN(n_5_923));
   NAND2_X1 i_5_1200 (.A1(n_5_842), .A2(n_5_387), .ZN(n_5_924));
   INV_X1 i_5_1201 (.A(n_5_3563), .ZN(n_5_925));
   INV_X1 i_5_1202 (.A(n_5_2568), .ZN(n_5_926));
   NAND2_X1 i_5_758 (.A1(n_5_925), .A2(n_5_926), .ZN(n_5_927));
   NAND3_X1 i_5_1204 (.A1(n_5_3784), .A2(n_5_717), .A3(n_5_4029), .ZN(n_5_928));
   NAND2_X1 i_5_1205 (.A1(n_5_745), .A2(n_5_3785), .ZN(n_5_929));
   NAND2_X1 i_5_1206 (.A1(n_5_928), .A2(n_5_929), .ZN(n_5_930));
   NAND2_X1 i_5_1207 (.A1(n_5_3776), .A2(n_5_674), .ZN(n_5_3141));
   NAND2_X1 i_5_1208 (.A1(n_5_740), .A2(m[6]), .ZN(n_5_931));
   INV_X1 i_5_1209 (.A(n_5_931), .ZN(n_5_932));
   NAND2_X1 i_5_1210 (.A1(n_5_4694), .A2(n_5_932), .ZN(n_5_933));
   INV_X1 i_5_1211 (.A(m[14]), .ZN(n_5_1806));
   INV_X1 i_5_1212 (.A(m[15]), .ZN(n_5_934));
   INV_X1 i_5_795 (.A(n_5_4155), .ZN(n_5_935));
   INV_X1 i_5_1214 (.A(m[10]), .ZN(n_5_936));
   INV_X1 i_5_1215 (.A(n_5_3377), .ZN(n_5_937));
   INV_X1 i_5_1216 (.A(m[13]), .ZN(n_5_938));
   NAND2_X1 i_5_1217 (.A1(n_5_3399), .A2(m[14]), .ZN(n_5_1817));
   INV_X1 i_5_1218 (.A(n_5_3399), .ZN(n_5_1819));
   INV_X1 i_5_1219 (.A(n_5_943), .ZN(n_5_939));
   INV_X1 i_5_1220 (.A(n_5_972), .ZN(n_5_1820));
   XNOR2_X1 i_5_1221 (.A(n_5_1002), .B(m[1]), .ZN(n_5_940));
   XNOR2_X1 i_5_1222 (.A(n_5_3365), .B(n_5_940), .ZN(n_5_3142));
   XNOR2_X1 i_5_1223 (.A(m[14]), .B(n_5_934), .ZN(n_5_3143));
   INV_X1 i_5_1224 (.A(m[14]), .ZN(n_5_941));
   INV_X1 i_5_1225 (.A(n_5_3399), .ZN(n_5_942));
   NAND2_X1 i_5_1226 (.A1(n_5_968), .A2(n_5_969), .ZN(n_5_943));
   AOI21_X1 i_5_1227 (.A(n_5_3751), .B1(n_5_976), .B2(n_5_944), .ZN(n_5_3355));
   INV_X1 i_5_1228 (.A(n_5_991), .ZN(n_5_944));
   AOI21_X1 i_5_1229 (.A(n_5_1002), .B1(n_5_3365), .B2(m[1]), .ZN(n_5_945));
   NAND2_X1 i_5_1230 (.A1(n_5_982), .A2(n_5_966), .ZN(n_5_3356));
   AOI21_X1 i_5_1231 (.A(n_5_973), .B1(n_5_995), .B2(n_5_993), .ZN(n_5_3357));
   OAI21_X1 i_5_797 (.A(n_5_971), .B1(n_5_977), .B2(n_5_957), .ZN(n_5_4057));
   XNOR2_X1 i_5_675 (.A(n_5_3067), .B(n_5_3080), .ZN(n_5_3147));
   XNOR2_X1 i_5_1234 (.A(n_5_946), .B(n_5_947), .ZN(n_5_3148));
   XNOR2_X1 i_5_1235 (.A(n_5_3377), .B(m[13]), .ZN(n_5_946));
   NAND2_X1 i_5_1236 (.A1(n_5_3088), .A2(n_5_3199), .ZN(n_5_947));
   NAND2_X1 i_5_1237 (.A1(n_5_951), .A2(n_5_948), .ZN(n_5_3149));
   OAI21_X1 i_5_1238 (.A(n_5_955), .B1(n_5_950), .B2(n_5_949), .ZN(n_5_948));
   NOR2_X1 i_5_1239 (.A1(n_5_3399), .A2(n_5_941), .ZN(n_5_949));
   INV_X1 i_5_1240 (.A(n_5_953), .ZN(n_5_950));
   NAND3_X1 i_5_1241 (.A1(n_5_954), .A2(n_5_953), .A3(n_5_952), .ZN(n_5_951));
   NAND2_X1 i_5_1242 (.A1(n_5_942), .A2(m[14]), .ZN(n_5_952));
   NAND2_X1 i_5_1243 (.A1(n_5_3399), .A2(n_5_941), .ZN(n_5_953));
   INV_X1 i_5_1244 (.A(n_5_955), .ZN(n_5_954));
   NAND2_X1 i_5_1245 (.A1(n_5_956), .A2(n_5_1844), .ZN(n_5_955));
   NAND3_X1 i_5_1246 (.A1(n_5_3088), .A2(n_5_972), .A3(n_5_3199), .ZN(n_5_956));
   NOR2_X1 i_5_1247 (.A1(n_5_3983), .A2(m[11]), .ZN(n_5_1826));
   AOI21_X1 i_5_1248 (.A(n_5_957), .B1(n_5_3983), .B2(m[11]), .ZN(n_5_1828));
   INV_X1 i_5_806 (.A(n_5_958), .ZN(n_5_957));
   NAND2_X1 i_5_811 (.A1(n_5_4155), .A2(m[10]), .ZN(n_5_958));
   NAND2_X1 i_5_790 (.A1(n_5_996), .A2(n_5_960), .ZN(n_5_959));
   OAI21_X1 i_5_809 (.A(n_5_995), .B1(n_5_973), .B2(n_5_961), .ZN(n_5_960));
   AOI21_X1 i_5_815 (.A(n_5_963), .B1(n_5_4145), .B2(n_5_962), .ZN(n_5_961));
   INV_X1 i_5_816 (.A(n_5_980), .ZN(n_5_962));
   INV_X1 i_5_817 (.A(n_5_4146), .ZN(n_5_963));
   NAND3_X1 i_5_818 (.A1(n_5_996), .A2(n_5_978), .A3(n_5_965), .ZN(n_5_964));
   AND3_X1 i_5_830 (.A1(n_5_994), .A2(n_5_4145), .A3(n_5_979), .ZN(n_5_965));
   NAND2_X1 i_5_1258 (.A1(n_5_3381), .A2(m[3]), .ZN(n_5_966));
   OAI22_X1 i_5_1259 (.A1(n_5_939), .A2(n_5_1000), .B1(n_5_969), .B2(n_5_968), 
      .ZN(n_5_967));
   INV_X1 i_5_1260 (.A(n_5_3365), .ZN(n_5_968));
   INV_X1 i_5_1261 (.A(m[1]), .ZN(n_5_969));
   INV_X1 i_5_837 (.A(n_5_4135), .ZN(n_5_970));
   NAND2_X1 i_5_855 (.A1(n_5_935), .A2(n_5_936), .ZN(n_5_971));
   NAND2_X1 i_5_1264 (.A1(n_5_3377), .A2(m[13]), .ZN(n_5_972));
   NAND2_X1 i_5_1265 (.A1(n_5_937), .A2(n_5_938), .ZN(n_5_1844));
   NOR2_X1 i_5_852 (.A1(n_5_4192), .A2(m[6]), .ZN(n_5_973));
   INV_X1 i_5_1267 (.A(m[6]), .ZN(n_5_974));
   INV_X1 i_5_1268 (.A(n_5_3751), .ZN(n_5_975));
   NAND2_X1 i_5_1269 (.A1(n_5_4101), .A2(m[2]), .ZN(n_5_976));
   INV_X1 i_5_1270 (.A(m[12]), .ZN(n_5_1850));
   NAND2_X1 i_5_1271 (.A1(n_5_977), .A2(n_5_971), .ZN(n_5_1863));
   AOI21_X1 i_5_856 (.A(n_5_3849), .B1(n_5_3844), .B2(n_5_989), .ZN(n_5_977));
   INV_X1 i_5_854 (.A(n_5_1005), .ZN(n_5_978));
   INV_X1 i_5_887 (.A(n_5_981), .ZN(n_5_979));
   NAND2_X1 i_5_888 (.A1(n_5_3401), .A2(m[4]), .ZN(n_5_980));
   NOR2_X1 i_5_1276 (.A1(n_5_3401), .A2(m[4]), .ZN(n_5_981));
   OR2_X1 i_5_1277 (.A1(n_5_3381), .A2(m[3]), .ZN(n_5_982));
   INV_X1 i_5_1278 (.A(m[4]), .ZN(n_5_983));
   XNOR2_X1 i_5_1279 (.A(n_5_3401), .B(n_5_983), .ZN(n_5_984));
   NAND2_X1 i_5_1280 (.A1(n_5_984), .A2(n_5_3575), .ZN(n_5_985));
   XNOR2_X1 i_5_1281 (.A(m[4]), .B(m[3]), .ZN(n_5_986));
   INV_X1 i_5_1282 (.A(n_5_3401), .ZN(n_5_987));
   XNOR2_X1 i_5_1283 (.A(n_5_1127), .B(n_5_987), .ZN(n_5_988));
   OAI21_X1 i_5_760 (.A(n_5_985), .B1(n_5_988), .B2(n_5_3575), .ZN(n_5_3151));
   NAND2_X1 i_5_913 (.A1(n_5_4108), .A2(m[9]), .ZN(n_5_989));
   AOI21_X1 i_5_1286 (.A(n_5_945), .B1(n_5_969), .B2(n_5_968), .ZN(n_5_990));
   XNOR2_X1 i_5_1287 (.A(n_5_3750), .B(n_5_990), .ZN(n_5_3152));
   AOI21_X1 i_5_1288 (.A(n_5_945), .B1(n_5_969), .B2(n_5_968), .ZN(n_5_991));
   INV_X1 i_5_1289 (.A(m[9]), .ZN(n_5_992));
   OAI21_X1 i_5_1290 (.A(n_5_4145), .B1(n_5_1004), .B2(n_5_963), .ZN(n_5_993));
   NAND2_X1 i_5_928 (.A1(n_5_3909), .A2(n_5_974), .ZN(n_5_994));
   NAND2_X1 i_5_937 (.A1(n_5_4192), .A2(m[6]), .ZN(n_5_995));
   INV_X1 i_5_1293 (.A(m[6]), .ZN(n_5_3359));
   INV_X1 i_5_1294 (.A(n_5_974), .ZN(n_5_1871));
   OR2_X1 i_5_941 (.A1(n_5_3372), .A2(m[7]), .ZN(n_5_996));
   NAND2_X1 i_5_942 (.A1(n_5_3372), .A2(m[7]), .ZN(n_5_997));
   XNOR2_X1 i_5_1297 (.A(n_5_3372), .B(m[7]), .ZN(n_5_3360));
   NAND2_X1 i_5_1298 (.A1(n_5_1871), .A2(n_5_3359), .ZN(n_5_998));
   INV_X1 i_5_1299 (.A(n_5_998), .ZN(n_5_999));
   OAI21_X1 i_5_1300 (.A(n_5_4145), .B1(n_5_1004), .B2(n_5_963), .ZN(n_5_2699));
   NAND2_X1 i_5_1301 (.A1(n_5_3364), .A2(m[0]), .ZN(n_5_1000));
   NAND2_X1 i_5_1302 (.A1(n_5_3364), .A2(m[0]), .ZN(n_5_1001));
   INV_X1 i_5_1303 (.A(n_5_1001), .ZN(n_5_1002));
   OAI21_X1 i_5_1304 (.A(n_5_980), .B1(n_5_3438), .B2(n_5_981), .ZN(n_5_1003));
   OAI21_X1 i_5_1305 (.A(n_5_980), .B1(n_5_3438), .B2(n_5_981), .ZN(n_5_1004));
   NAND2_X1 i_5_947 (.A1(n_5_982), .A2(n_5_3439), .ZN(n_5_1005));
   INV_X1 i_5_1307 (.A(n_5_999), .ZN(n_5_1923));
   NAND2_X1 i_5_1308 (.A1(n_5_975), .A2(n_5_967), .ZN(n_5_1007));
   NAND2_X1 i_5_1309 (.A1(n_5_975), .A2(n_5_967), .ZN(n_5_1008));
   NAND2_X1 i_5_1310 (.A1(n_5_2016), .A2(n_5_1036), .ZN(n_5_1009));
   NAND2_X1 i_5_1311 (.A1(n_5_1107), .A2(n_5_1038), .ZN(n_5_1010));
   NAND2_X1 i_5_1312 (.A1(n_5_3063), .A2(n_5_1039), .ZN(n_5_1011));
   NAND3_X1 i_5_1313 (.A1(n_5_1009), .A2(n_5_1010), .A3(n_5_1011), .ZN(n_5_3364));
   NAND2_X1 i_5_1314 (.A1(n_5_2028), .A2(n_5_1036), .ZN(n_5_1012));
   NAND2_X1 i_5_1315 (.A1(n_5_3140), .A2(n_5_1039), .ZN(n_5_1013));
   NAND3_X1 i_5_1316 (.A1(n_5_3235), .A2(n_5_1012), .A3(n_5_1013), .ZN(n_5_3365));
   NAND2_X1 i_5_1317 (.A1(n_5_2024), .A2(n_5_1036), .ZN(n_5_3366));
   NAND2_X1 i_5_1318 (.A1(n_5_3398), .A2(n_5_1039), .ZN(n_5_3367));
   NAND2_X1 i_5_1319 (.A1(n_5_1962), .A2(n_5_1036), .ZN(n_5_1014));
   NAND2_X1 i_5_1320 (.A1(n_5_3068), .A2(n_5_1039), .ZN(n_5_1015));
   NAND2_X1 i_5_1321 (.A1(n_5_3746), .A2(n_5_1039), .ZN(n_5_1924));
   NAND2_X1 i_5_957 (.A1(n_5_1976), .A2(n_5_1036), .ZN(n_5_1016));
   NAND2_X1 i_5_958 (.A1(n_5_1049), .A2(n_5_1038), .ZN(n_5_1017));
   NAND2_X1 i_5_1324 (.A1(n_5_3418), .A2(n_5_1039), .ZN(n_5_1018));
   NAND2_X1 i_5_959 (.A1(n_5_2008), .A2(n_5_1036), .ZN(n_5_1019));
   NAND2_X1 i_5_972 (.A1(n_5_1051), .A2(n_5_1038), .ZN(n_5_1020));
   NAND2_X1 i_5_1327 (.A1(n_5_4394), .A2(n_5_1039), .ZN(n_5_1021));
   NAND2_X1 i_5_1025 (.A1(n_5_1978), .A2(n_5_1036), .ZN(n_5_1022));
   NAND2_X1 i_5_1329 (.A1(n_5_3291), .A2(n_5_1039), .ZN(n_5_1023));
   NAND3_X1 i_5_1065 (.A1(n_5_3046), .A2(n_5_1022), .A3(n_5_1023), .ZN(n_5_3372));
   NAND2_X1 i_5_1331 (.A1(n_5_1052), .A2(n_5_1038), .ZN(n_5_1024));
   NAND2_X1 i_5_1332 (.A1(n_5_1981), .A2(n_5_1036), .ZN(n_5_1025));
   NAND2_X1 i_5_1333 (.A1(n_5_3406), .A2(n_5_1039), .ZN(n_5_1026));
   NAND2_X1 i_5_1066 (.A1(n_5_1053), .A2(n_5_1038), .ZN(n_5_1027));
   NAND2_X1 i_5_1335 (.A1(n_5_3382), .A2(n_5_1039), .ZN(n_5_1028));
   NAND2_X1 i_5_1067 (.A1(n_5_1058), .A2(n_5_1038), .ZN(n_5_1029));
   NAND2_X1 i_5_1337 (.A1(n_5_3229), .A2(n_5_1039), .ZN(n_5_1030));
   NAND2_X1 i_5_945 (.A1(n_5_1062), .A2(n_5_1038), .ZN(n_5_456));
   NAND2_X1 i_5_1094 (.A1(n_5_3320), .A2(n_5_1039), .ZN(n_5_460));
   NAND2_X1 i_5_1233 (.A1(n_5_1096), .A2(n_5_1038), .ZN(n_5_4059));
   NAND2_X1 i_5_1272 (.A1(n_5_1996), .A2(n_5_1036), .ZN(n_5_4060));
   NAND2_X1 i_5_1343 (.A1(n_5_3219), .A2(n_5_1039), .ZN(n_5_4061));
   NAND2_X1 i_5_1344 (.A1(n_5_1069), .A2(n_5_1038), .ZN(n_5_1033));
   NAND2_X1 i_5_1345 (.A1(n_5_1997), .A2(n_5_1036), .ZN(n_5_1034));
   NAND3_X1 i_5_1346 (.A1(n_5_1033), .A2(n_5_1034), .A3(n_5_1938), .ZN(n_5_3377));
   INV_X1 i_5_1347 (.A(r[4]), .ZN(n_5_1035));
   NOR2_X1 i_5_1348 (.A1(r[5]), .A2(n_5_1035), .ZN(n_5_1036));
   NAND2_X1 i_5_1349 (.A1(r[5]), .A2(n_5_1035), .ZN(n_5_1037));
   INV_X1 i_5_1350 (.A(n_5_1037), .ZN(n_5_1038));
   XNOR2_X1 i_5_1351 (.A(r[5]), .B(r[4]), .ZN(n_5_1039));
   NAND2_X1 i_5_1352 (.A1(n_5_2167), .A2(n_5_1039), .ZN(n_5_1938));
   INV_X1 i_5_1353 (.A(n_53), .ZN(n_5_1040));
   INV_X1 i_5_1354 (.A(n_54), .ZN(n_5_1041));
   INV_X1 i_5_1355 (.A(n_5_3746), .ZN(n_5_1042));
   INV_X1 i_5_1356 (.A(n_66), .ZN(n_5_1043));
   INV_X1 i_5_1357 (.A(n_75), .ZN(n_5_1044));
   INV_X1 i_5_1358 (.A(n_61), .ZN(n_5_1045));
   INV_X1 i_5_1359 (.A(n_5_2167), .ZN(n_5_1046));
   NAND2_X1 i_5_1360 (.A1(n_5_3304), .A2(n_5_1953), .ZN(n_5_1047));
   AOI21_X1 i_5_1102 (.A(n_5_1104), .B1(n_5_1047), .B2(n_5_3265), .ZN(n_5_1048));
   XNOR2_X1 i_5_1104 (.A(n_5_1048), .B(n_5_1091), .ZN(n_5_1049));
   NAND2_X1 i_5_1363 (.A1(n_5_3284), .A2(n_5_3330), .ZN(n_5_1050));
   XNOR2_X1 i_5_1364 (.A(n_5_1087), .B(n_5_1050), .ZN(n_5_1051));
   INV_X1 i_5_1098 (.A(n_5_1086), .ZN(n_5_4062));
   NAND2_X1 i_5_1099 (.A1(n_5_3284), .A2(n_5_3573), .ZN(n_5_4063));
   XOR2_X1 i_5_1367 (.A(n_5_3404), .B(n_5_1110), .Z(n_5_1052));
   XNOR2_X1 i_5_1368 (.A(n_5_1090), .B(n_5_1112), .ZN(n_5_1053));
   INV_X1 i_5_1369 (.A(n_5_3038), .ZN(n_5_1054));
   NOR2_X1 i_5_1101 (.A1(n_5_3229), .A2(n_76), .ZN(n_5_1055));
   NOR2_X1 i_5_1371 (.A1(n_5_1054), .A2(n_5_1055), .ZN(n_5_1056));
   NAND2_X1 i_5_1372 (.A1(n_5_1085), .A2(n_5_1088), .ZN(n_5_1057));
   XNOR2_X1 i_5_1373 (.A(n_5_1056), .B(n_5_1057), .ZN(n_5_1058));
   INV_X1 i_5_1115 (.A(n_5_1089), .ZN(n_5_1059));
   AOI21_X1 i_5_1118 (.A(n_5_1059), .B1(n_5_1088), .B2(n_5_1113), .ZN(n_5_1060));
   OAI21_X1 i_5_1186 (.A(n_5_3038), .B1(n_5_1060), .B2(n_5_1055), .ZN(n_5_1061));
   XNOR2_X1 i_5_1213 (.A(n_5_3319), .B(n_5_1061), .ZN(n_5_1062));
   XNOR2_X1 i_5_1092 (.A(n_5_3219), .B(n_61), .ZN(n_5_1063));
   NAND2_X1 i_5_1379 (.A1(n_5_3318), .A2(n_5_1044), .ZN(n_5_1064));
   XNOR2_X1 i_5_1380 (.A(n_5_2167), .B(n_53), .ZN(n_5_1065));
   NAND2_X1 i_5_1381 (.A1(n_5_3219), .A2(n_61), .ZN(n_5_1066));
   NAND3_X1 i_5_1382 (.A1(n_5_1065), .A2(n_5_1108), .A3(n_5_1095), .ZN(n_5_1067));
   AND2_X1 i_5_1383 (.A1(n_5_1095), .A2(n_5_1108), .ZN(n_5_1068));
   OAI21_X1 i_5_1384 (.A(n_5_1067), .B1(n_5_1068), .B2(n_5_1065), .ZN(n_5_1069));
   XOR2_X1 i_5_1385 (.A(n_5_1041), .B(n_53), .Z(n_5_1070));
   INV_X1 i_5_1386 (.A(n_5_1066), .ZN(n_5_1071));
   AOI21_X1 i_5_1387 (.A(n_5_1071), .B1(n_5_1040), .B2(n_5_1046), .ZN(n_5_1072));
   OAI21_X1 i_5_1388 (.A(n_5_1072), .B1(n_5_1097), .B2(n_5_1117), .ZN(n_5_1073));
   OAI21_X1 i_5_1389 (.A(n_5_1070), .B1(n_5_1098), .B2(n_5_1099), .ZN(n_5_3157));
   NAND2_X1 i_5_1390 (.A1(n_5_3140), .A2(n_5_3329), .ZN(n_5_1074));
   INV_X1 i_5_1391 (.A(n_5_3329), .ZN(n_5_1942));
   NAND2_X1 i_5_1392 (.A1(n_5_1944), .A2(n_5_1953), .ZN(n_5_1075));
   NOR2_X1 i_5_1232 (.A1(n_5_3520), .A2(n_5_1075), .ZN(n_5_4064));
   INV_X1 i_5_1249 (.A(n_5_3286), .ZN(n_5_1076));
   NAND2_X1 i_5_1395 (.A1(n_5_1093), .A2(n_5_1101), .ZN(n_5_1943));
   NAND2_X1 i_5_1250 (.A1(n_5_3406), .A2(n_55), .ZN(n_5_1077));
   NOR2_X1 i_5_1285 (.A1(n_5_3406), .A2(n_55), .ZN(n_5_1078));
   OAI21_X1 i_5_1398 (.A(n_5_1119), .B1(n_5_3406), .B2(n_55), .ZN(n_5_1079));
   INV_X1 i_5_1399 (.A(n_55), .ZN(n_5_1080));
   NOR2_X1 i_5_1400 (.A1(n_5_3450), .A2(n_5_1080), .ZN(n_5_1081));
   NAND2_X1 i_5_1401 (.A1(n_5_3450), .A2(n_5_1080), .ZN(n_5_1082));
   AOI21_X1 i_5_1402 (.A(n_5_1081), .B1(n_5_3406), .B2(n_5_1082), .ZN(n_5_1083));
   NAND2_X1 i_5_1403 (.A1(n_5_3382), .A2(n_73), .ZN(n_5_1084));
   NAND3_X1 i_5_1404 (.A1(n_5_1079), .A2(n_5_1083), .A3(n_5_1084), .ZN(n_5_1085));
   NAND2_X1 i_5_1405 (.A1(n_5_4394), .A2(n_69), .ZN(n_5_1086));
   XNOR2_X1 i_5_1406 (.A(n_5_4394), .B(n_69), .ZN(n_5_1087));
   OR2_X1 i_5_1338 (.A1(n_5_3382), .A2(n_73), .ZN(n_5_1088));
   NAND2_X1 i_5_1339 (.A1(n_5_3382), .A2(n_73), .ZN(n_5_1089));
   XNOR2_X1 i_5_1409 (.A(n_5_3382), .B(n_73), .ZN(n_5_1090));
   NAND2_X1 i_5_1107 (.A1(n_5_3518), .A2(n_5_3264), .ZN(n_5_1091));
   INV_X1 i_5_1411 (.A(n_5_2568), .ZN(n_5_1092));
   NAND2_X1 i_5_1412 (.A1(n_5_3059), .A2(n_5_1092), .ZN(n_5_1093));
   AOI22_X1 i_5_1413 (.A1(n_5_1061), .A2(n_5_1064), .B1(n_5_3320), .B2(n_75), 
      .ZN(n_5_1094));
   NAND2_X1 i_5_1414 (.A1(n_5_1066), .A2(n_5_1094), .ZN(n_5_1095));
   XOR2_X1 i_5_1394 (.A(n_5_1063), .B(n_5_1097), .Z(n_5_1096));
   AOI22_X1 i_5_1341 (.A1(n_5_1061), .A2(n_5_1064), .B1(n_5_3320), .B2(n_75), 
      .ZN(n_5_1097));
   INV_X1 i_5_1417 (.A(n_5_1073), .ZN(n_5_1098));
   AND2_X1 i_5_1418 (.A1(n_5_2167), .A2(n_53), .ZN(n_5_1099));
   AOI21_X1 i_5_1419 (.A(n_5_1070), .B1(n_5_2167), .B2(n_53), .ZN(n_5_1100));
   NAND2_X1 i_5_1420 (.A1(n_5_1073), .A2(n_5_1100), .ZN(n_5_3158));
   INV_X1 i_5_1421 (.A(n_5_1105), .ZN(n_5_1101));
   INV_X1 i_5_1422 (.A(n_5_2568), .ZN(n_5_1102));
   NAND2_X1 i_5_1423 (.A1(n_5_1042), .A2(n_5_1043), .ZN(n_5_1944));
   NAND2_X1 i_5_1424 (.A1(n_5_1042), .A2(n_5_1043), .ZN(n_5_1103));
   INV_X1 i_5_1425 (.A(n_5_1103), .ZN(n_5_1104));
   BUF_X1 i_5_1426 (.A(n_5_3425), .Z(n_5_1105));
   XNOR2_X1 i_5_1427 (.A(n_5_3425), .B(n_5_1102), .ZN(n_5_1106));
   XNOR2_X1 i_5_1428 (.A(n_5_1106), .B(n_5_3063), .ZN(n_5_1107));
   NAND2_X1 i_5_1429 (.A1(n_5_1115), .A2(n_5_1045), .ZN(n_5_1108));
   INV_X1 i_5_1430 (.A(n_5_4062), .ZN(n_5_1109));
   NAND2_X1 i_5_1431 (.A1(n_5_1121), .A2(n_5_1109), .ZN(n_5_1945));
   OAI21_X1 i_5_1432 (.A(n_5_1076), .B1(n_5_4337), .B2(n_5_3452), .ZN(n_5_1110));
   OR2_X1 i_5_1433 (.A1(n_5_3068), .A2(n_58), .ZN(n_5_1953));
   XNOR2_X1 i_5_1434 (.A(n_5_3068), .B(n_58), .ZN(n_5_3379));
   NAND2_X1 i_5_1435 (.A1(n_5_3422), .A2(n_5_3423), .ZN(n_5_3380));
   AOI21_X1 i_5_1436 (.A(n_5_3452), .B1(n_5_4337), .B2(n_5_1076), .ZN(n_5_1111));
   AOI21_X1 i_5_1437 (.A(n_5_1078), .B1(n_5_1111), .B2(n_5_1077), .ZN(n_5_1112));
   OAI21_X1 i_5_1340 (.A(n_5_1077), .B1(n_5_1114), .B2(n_5_1078), .ZN(n_5_1113));
   AOI21_X1 i_5_1362 (.A(n_5_3452), .B1(n_5_4337), .B2(n_5_1076), .ZN(n_5_1114));
   INV_X1 i_5_1440 (.A(n_5_3219), .ZN(n_5_1115));
   INV_X1 i_5_1441 (.A(n_5_1045), .ZN(n_5_1116));
   NOR2_X1 i_5_1442 (.A1(n_5_3219), .A2(n_5_1116), .ZN(n_5_1117));
   NOR2_X1 i_5_1443 (.A1(n_5_3291), .A2(n_60), .ZN(n_5_1118));
   OAI22_X1 i_5_1444 (.A1(n_5_4333), .A2(n_5_1118), .B1(n_5_1118), .B2(n_5_4334), 
      .ZN(n_5_1119));
   OR2_X1 i_5_1445 (.A1(n_5_4394), .A2(n_69), .ZN(n_5_1120));
   OAI21_X1 i_5_1446 (.A(n_5_1120), .B1(n_5_4063), .B2(n_5_4064), .ZN(n_5_1121));
   OAI21_X1 i_5_1447 (.A(n_5_3058), .B1(n_5_3056), .B2(n_5_3425), .ZN(n_5_1956));
   NAND3_X1 i_5_1448 (.A1(n_5_1019), .A2(n_5_1020), .A3(n_5_1021), .ZN(n_5_1122));
   INV_X1 i_5_1449 (.A(n_5_1122), .ZN(n_5_1960));
   NAND3_X1 i_5_1450 (.A1(n_5_3766), .A2(n_5_1014), .A3(n_5_1015), .ZN(n_5_3381));
   NAND3_X1 i_5_1451 (.A1(n_5_3766), .A2(n_5_1014), .A3(n_5_1015), .ZN(n_5_1123));
   INV_X1 i_5_1452 (.A(n_5_1123), .ZN(n_5_1124));
   NAND2_X1 i_5_1453 (.A1(n_5_1124), .A2(n_5_986), .ZN(n_5_1125));
   NAND2_X1 i_5_1454 (.A1(n_5_1123), .A2(m[4]), .ZN(n_5_1126));
   NAND2_X1 i_5_1455 (.A1(n_5_1125), .A2(n_5_1126), .ZN(n_5_1127));
   XNOR2_X1 i_5_1456 (.A(n_5_3844), .B(n_5_3850), .ZN(n_5_3160));
   AOI21_X1 i_5_1129 (.A(n_5_3849), .B1(n_5_3845), .B2(n_5_989), .ZN(n_5_3864));
   XNOR2_X1 i_5_1458 (.A(n_5_3071), .B(n_5_3411), .ZN(n_5_1128));
   NAND2_X1 i_5_1459 (.A1(n_5_1128), .A2(n_5_1038), .ZN(n_5_3383));
   XNOR2_X1 i_5_1460 (.A(n_5_1129), .B(n_5_1189), .ZN(n_5_1962));
   NAND2_X1 i_5_1461 (.A1(n_5_3043), .A2(n_5_3460), .ZN(n_5_1129));
   XOR2_X1 i_5_1462 (.A(n_5_3036), .B(n_5_3254), .Z(n_5_1968));
   XOR2_X1 i_5_1162 (.A(n_5_3373), .B(n_5_1143), .Z(n_5_1976));
   XNOR2_X1 i_5_1464 (.A(n_5_3290), .B(n_5_1203), .ZN(n_5_1978));
   XOR2_X1 i_5_1465 (.A(n_5_1204), .B(n_5_3405), .Z(n_5_1981));
   NAND2_X1 i_5_1466 (.A1(n_5_3233), .A2(n_5_2972), .ZN(n_5_1130));
   XNOR2_X1 i_5_1407 (.A(n_5_1131), .B(n_5_1164), .ZN(n_5_1996));
   NAND2_X1 i_5_1468 (.A1(n_5_1149), .A2(n_5_2949), .ZN(n_5_1131));
   XNOR2_X1 i_5_1469 (.A(n_5_1132), .B(n_5_1172), .ZN(n_5_1997));
   OAI21_X1 i_5_1470 (.A(n_5_1149), .B1(n_5_1164), .B2(n_5_2951), .ZN(n_5_1132));
   NAND2_X1 i_5_1471 (.A1(n_5_1133), .A2(n_5_1135), .ZN(n_5_1998));
   NAND2_X1 i_5_1472 (.A1(n_5_1134), .A2(n_5_1137), .ZN(n_5_1133));
   NAND2_X1 i_5_1473 (.A1(n_5_1192), .A2(n_5_1170), .ZN(n_5_1134));
   NAND3_X1 i_5_1474 (.A1(n_5_1192), .A2(n_5_1170), .A3(n_5_1136), .ZN(n_5_1135));
   INV_X1 i_5_1475 (.A(n_5_1137), .ZN(n_5_1136));
   XNOR2_X1 i_5_1476 (.A(n_5_1138), .B(m[14]), .ZN(n_5_1137));
   INV_X1 i_5_1477 (.A(m[15]), .ZN(n_5_1138));
   INV_X1 i_5_1478 (.A(m[12]), .ZN(n_5_1139));
   OAI21_X1 i_5_1365 (.A(n_5_3233), .B1(n_5_1141), .B2(n_5_1148), .ZN(n_5_1140));
   AOI21_X1 i_5_1480 (.A(n_5_1153), .B1(n_5_1142), .B2(n_5_1199), .ZN(n_5_1141));
   NAND2_X1 i_5_1481 (.A1(n_5_1207), .A2(n_5_1155), .ZN(n_5_1142));
   NAND2_X1 i_5_1163 (.A1(n_5_1144), .A2(n_5_1173), .ZN(n_5_1143));
   NAND2_X1 i_5_1180 (.A1(n_5_3254), .A2(n_5_1174), .ZN(n_5_1144));
   NAND2_X1 i_5_1484 (.A1(n_5_1211), .A2(m[0]), .ZN(n_5_1145));
   INV_X1 i_5_1485 (.A(n_5_1187), .ZN(n_5_1146));
   INV_X1 i_5_1486 (.A(n_5_3288), .ZN(n_5_1147));
   INV_X1 i_5_1487 (.A(n_5_2972), .ZN(n_5_1148));
   NAND2_X1 i_5_1488 (.A1(n_5_1150), .A2(n_5_1151), .ZN(n_5_1149));
   INV_X1 i_5_1489 (.A(n_5_3219), .ZN(n_5_1150));
   INV_X1 i_5_1490 (.A(m[13]), .ZN(n_5_1151));
   INV_X1 i_5_1491 (.A(m[3]), .ZN(n_5_1152));
   NOR2_X1 i_5_1492 (.A1(n_5_3382), .A2(m[10]), .ZN(n_5_1153));
   INV_X1 i_5_1493 (.A(m[10]), .ZN(n_5_1154));
   INV_X1 i_5_1494 (.A(m[3]), .ZN(n_5_1999));
   INV_X1 i_5_1495 (.A(n_5_1152), .ZN(n_5_2005));
   OR2_X1 i_5_1496 (.A1(n_5_3406), .A2(m[9]), .ZN(n_5_1155));
   INV_X1 i_5_1497 (.A(m[1]), .ZN(n_5_1156));
   NAND2_X1 i_5_1498 (.A1(n_5_3060), .A2(n_5_1156), .ZN(n_5_1157));
   NAND2_X1 i_5_1499 (.A1(n_5_4394), .A2(m[7]), .ZN(n_5_1158));
   AOI21_X1 i_5_1500 (.A(n_5_4171), .B1(m[12]), .B2(n_5_3320), .ZN(n_5_1159));
   INV_X1 i_5_1501 (.A(n_5_3320), .ZN(n_5_1160));
   NAND2_X1 i_5_1502 (.A1(n_5_3320), .A2(m[12]), .ZN(n_5_1161));
   INV_X1 i_5_1503 (.A(n_5_1139), .ZN(n_5_1162));
   NOR2_X1 i_5_1504 (.A1(n_5_3320), .A2(n_5_1162), .ZN(n_5_1163));
   OAI21_X1 i_5_1505 (.A(n_5_1161), .B1(n_5_1140), .B2(n_5_1163), .ZN(n_5_1164));
   INV_X1 i_5_1506 (.A(m[7]), .ZN(n_5_1165));
   XNOR2_X1 i_5_1507 (.A(n_5_4394), .B(n_5_1165), .ZN(n_5_1166));
   INV_X1 i_5_1508 (.A(n_5_3476), .ZN(n_5_1167));
   NAND2_X1 i_5_1509 (.A1(n_5_1166), .A2(n_5_1167), .ZN(n_5_1168));
   XNOR2_X1 i_5_1510 (.A(n_5_1193), .B(n_5_4394), .ZN(n_5_1169));
   OAI21_X1 i_5_1511 (.A(n_5_1168), .B1(n_5_1169), .B2(n_5_1167), .ZN(n_5_2008));
   OR2_X1 i_5_1512 (.A1(m[14]), .A2(n_5_2167), .ZN(n_5_1170));
   INV_X1 i_5_1513 (.A(m[14]), .ZN(n_5_1171));
   XNOR2_X1 i_5_1514 (.A(n_5_2167), .B(n_5_1171), .ZN(n_5_1172));
   OR2_X1 i_5_1181 (.A1(n_5_3746), .A2(m[5]), .ZN(n_5_1173));
   NAND2_X1 i_5_1189 (.A1(n_5_3746), .A2(m[5]), .ZN(n_5_1174));
   NAND2_X1 i_5_1517 (.A1(n_5_2167), .A2(m[14]), .ZN(n_5_1175));
   INV_X1 i_5_1518 (.A(n_5_1175), .ZN(n_5_1176));
   NAND2_X1 i_5_1519 (.A1(n_5_1150), .A2(n_5_1151), .ZN(n_5_1177));
   INV_X1 i_5_1520 (.A(n_5_2949), .ZN(n_5_1178));
   NAND2_X1 i_5_1521 (.A1(n_5_1160), .A2(n_5_1139), .ZN(n_5_1179));
   OAI21_X1 i_5_1522 (.A(n_5_1177), .B1(n_5_1178), .B2(n_5_1179), .ZN(n_5_1180));
   NAND2_X1 i_5_1523 (.A1(n_5_2949), .A2(n_5_1149), .ZN(n_5_1181));
   INV_X1 i_5_1524 (.A(n_5_1181), .ZN(n_5_1182));
   INV_X1 i_5_1525 (.A(n_5_1157), .ZN(n_5_1183));
   INV_X1 i_5_1526 (.A(n_5_1145), .ZN(n_5_1184));
   NAND2_X1 i_5_1527 (.A1(n_5_1183), .A2(n_5_1184), .ZN(n_5_1185));
   OAI21_X1 i_5_1528 (.A(n_5_1185), .B1(n_5_1200), .B2(n_5_1183), .ZN(n_5_2016));
   OR2_X1 i_5_1529 (.A1(n_5_3140), .A2(m[2]), .ZN(n_5_1186));
   NAND2_X1 i_5_1530 (.A1(n_5_3140), .A2(m[2]), .ZN(n_5_1187));
   XNOR2_X1 i_5_1531 (.A(n_5_3140), .B(m[2]), .ZN(n_5_1188));
   AOI21_X1 i_5_1532 (.A(n_5_3075), .B1(n_5_3076), .B2(n_5_2029), .ZN(n_5_1189));
   NAND2_X1 i_5_1533 (.A1(n_5_1182), .A2(n_5_1159), .ZN(n_5_1190));
   NOR2_X1 i_5_1534 (.A1(n_5_1180), .A2(n_5_1176), .ZN(n_5_1191));
   NAND2_X1 i_5_1535 (.A1(n_5_1190), .A2(n_5_1191), .ZN(n_5_1192));
   XNOR2_X1 i_5_1536 (.A(n_5_2933), .B(n_5_1165), .ZN(n_5_1193));
   NAND2_X1 i_5_1537 (.A1(n_5_2005), .A2(n_5_1999), .ZN(n_5_1194));
   INV_X1 i_5_1538 (.A(n_5_1194), .ZN(n_5_2023));
   NAND2_X1 i_5_1539 (.A1(n_5_3073), .A2(n_5_3074), .ZN(n_5_1195));
   OAI21_X1 i_5_1540 (.A(n_5_1186), .B1(n_5_1198), .B2(n_5_1146), .ZN(n_5_1196));
   XNOR2_X1 i_5_1541 (.A(n_5_1195), .B(n_5_1196), .ZN(n_5_2024));
   AOI21_X1 i_5_1542 (.A(n_5_3061), .B1(n_5_1201), .B2(n_5_1145), .ZN(n_5_1197));
   XNOR2_X1 i_5_1543 (.A(n_5_1188), .B(n_5_1198), .ZN(n_5_2028));
   OAI21_X1 i_5_1544 (.A(n_5_1186), .B1(n_5_1146), .B2(n_5_1197), .ZN(n_5_2029));
   AOI21_X1 i_5_1545 (.A(n_5_3061), .B1(n_5_1201), .B2(n_5_1145), .ZN(n_5_1198));
   NAND2_X1 i_5_1546 (.A1(n_5_3382), .A2(m[10]), .ZN(n_5_1199));
   INV_X1 i_5_1547 (.A(m[10]), .ZN(n_5_2031));
   INV_X1 i_5_1548 (.A(n_5_1154), .ZN(n_5_2032));
   XNOR2_X1 i_5_1549 (.A(n_5_3062), .B(n_5_1184), .ZN(n_5_1200));
   NAND2_X1 i_5_1550 (.A1(n_5_3063), .A2(m[1]), .ZN(n_5_1201));
   NOR2_X1 i_5_1551 (.A1(n_5_4394), .A2(m[7]), .ZN(n_5_1202));
   OAI22_X1 i_5_1552 (.A1(n_5_3475), .A2(n_5_1202), .B1(n_5_1158), .B2(n_5_1202), 
      .ZN(n_5_1203));
   OAI21_X1 i_5_1553 (.A(n_5_3289), .B1(n_5_1203), .B2(n_5_1147), .ZN(n_5_1204));
   OAI21_X1 i_5_1554 (.A(n_5_3289), .B1(n_5_1147), .B2(n_5_1203), .ZN(n_5_1205));
   NAND2_X1 i_5_1555 (.A1(n_5_3406), .A2(m[9]), .ZN(n_5_1206));
   NAND2_X1 i_5_1556 (.A1(n_5_1205), .A2(n_5_1206), .ZN(n_5_1207));
   NAND2_X1 i_5_1557 (.A1(n_5_1946), .A2(n_5_3386), .ZN(n_5_1208));
   NAND2_X1 i_5_1558 (.A1(n_5_1973), .A2(n_5_3385), .ZN(n_5_1209));
   NAND2_X1 i_5_1559 (.A1(n_5_2006), .A2(n_5_2165), .ZN(n_5_1210));
   NAND3_X1 i_5_1560 (.A1(n_5_1208), .A2(n_5_1209), .A3(n_5_1210), .ZN(n_5_1211));
   NAND2_X1 i_5_1561 (.A1(n_5_1947), .A2(n_5_3386), .ZN(n_5_2049));
   NAND2_X1 i_5_1562 (.A1(n_5_1974), .A2(n_5_3385), .ZN(n_5_2050));
   NAND2_X1 i_5_1563 (.A1(n_5_2002), .A2(n_5_2165), .ZN(n_5_2051));
   NAND2_X1 i_5_1564 (.A1(n_5_1980), .A2(n_5_3385), .ZN(n_5_2088));
   NAND2_X1 i_5_1565 (.A1(n_5_2012), .A2(n_5_2165), .ZN(n_5_2089));
   NAND2_X1 i_5_1566 (.A1(n_5_1987), .A2(n_5_3385), .ZN(n_5_2090));
   NAND2_X1 i_5_1567 (.A1(n_5_1719), .A2(n_5_2165), .ZN(n_5_2110));
   NAND2_X1 i_5_1568 (.A1(n_5_1784), .A2(n_5_2165), .ZN(n_5_1212));
   NAND2_X1 i_5_1569 (.A1(n_5_3029), .A2(n_5_2165), .ZN(n_5_3384));
   NAND2_X1 i_5_1251 (.A1(n_5_1984), .A2(n_5_3385), .ZN(n_5_1213));
   NAND2_X1 i_5_1252 (.A1(n_5_3113), .A2(n_5_2165), .ZN(n_5_2116));
   NAND2_X1 i_5_1572 (.A1(n_5_3168), .A2(n_5_2165), .ZN(n_5_2153));
   NAND2_X1 i_5_1366 (.A1(n_5_1952), .A2(n_5_3386), .ZN(n_5_2154));
   NAND2_X1 i_5_1574 (.A1(n_5_3297), .A2(n_5_2165), .ZN(n_5_2155));
   NAND2_X1 i_5_1575 (.A1(n_5_3816), .A2(n_5_3386), .ZN(n_5_2156));
   NAND2_X1 i_5_1576 (.A1(n_5_2007), .A2(n_5_3385), .ZN(n_5_2157));
   NAND2_X1 i_5_1577 (.A1(n_5_1751), .A2(n_5_2165), .ZN(n_5_2158));
   NAND2_X1 i_5_1578 (.A1(n_5_2013), .A2(n_5_2165), .ZN(n_5_2159));
   NAND2_X1 i_5_1370 (.A1(n_5_1954), .A2(n_5_3386), .ZN(n_5_2160));
   NAND2_X1 i_5_1374 (.A1(n_5_1977), .A2(n_5_3385), .ZN(n_5_2161));
   NAND2_X1 i_5_1581 (.A1(n_5_2017), .A2(n_5_2165), .ZN(n_5_2162));
   INV_X1 i_5_1582 (.A(r[3]), .ZN(n_5_1214));
   NOR2_X1 i_5_1583 (.A1(r[4]), .A2(n_5_1214), .ZN(n_5_3385));
   NAND2_X1 i_5_1584 (.A1(n_5_2984), .A2(n_5_3385), .ZN(n_5_1215));
   NAND2_X1 i_5_1585 (.A1(r[4]), .A2(n_5_1214), .ZN(n_5_1216));
   INV_X1 i_5_1586 (.A(n_5_1216), .ZN(n_5_3386));
   NAND2_X1 i_5_1587 (.A1(n_5_1958), .A2(n_5_3386), .ZN(n_5_1217));
   XNOR2_X1 i_5_1588 (.A(r[4]), .B(r[3]), .ZN(n_5_2165));
   NAND2_X1 i_5_1589 (.A1(n_5_464), .A2(n_5_2165), .ZN(n_5_2166));
   NAND3_X1 i_5_1590 (.A1(n_5_1215), .A2(n_5_1217), .A3(n_5_2166), .ZN(n_5_2167));
   INV_X1 i_5_1591 (.A(n_53), .ZN(n_5_1218));
   INV_X1 i_5_1592 (.A(n_54), .ZN(n_5_1219));
   INV_X1 i_5_1593 (.A(n_73), .ZN(n_5_1220));
   INV_X1 i_5_1594 (.A(n_5_2017), .ZN(n_5_1221));
   INV_X1 i_5_1595 (.A(n_61), .ZN(n_5_1222));
   INV_X1 i_5_1596 (.A(n_5_464), .ZN(n_5_1223));
   XNOR2_X1 i_5_1597 (.A(n_5_2006), .B(n_5_2568), .ZN(n_5_1224));
   XNOR2_X1 i_5_1598 (.A(n_5_3184), .B(n_5_1224), .ZN(n_5_1946));
   NAND2_X1 i_5_1599 (.A1(n_5_1226), .A2(n_5_1249), .ZN(n_5_1225));
   NAND2_X1 i_5_1600 (.A1(n_5_1223), .A2(n_5_1218), .ZN(n_5_1226));
   INV_X1 i_5_1601 (.A(n_53), .ZN(n_5_1227));
   NAND2_X1 i_5_1602 (.A1(n_5_1429), .A2(m[0]), .ZN(n_5_1228));
   NAND2_X1 i_5_1603 (.A1(n_5_2006), .A2(n_5_2568), .ZN(n_5_1229));
   INV_X1 i_5_1604 (.A(n_5_2006), .ZN(n_5_1230));
   INV_X1 i_5_1605 (.A(n_5_2568), .ZN(n_5_1231));
   AOI22_X1 i_5_1606 (.A1(n_5_1228), .A2(n_5_1229), .B1(n_5_1230), .B2(n_5_1231), 
      .ZN(n_5_1232));
   XNOR2_X1 i_5_1607 (.A(n_5_1290), .B(n_5_1232), .ZN(n_5_1947));
   NAND2_X1 i_5_1253 (.A1(n_5_1261), .A2(n_5_1260), .ZN(n_5_1950));
   AOI21_X1 i_5_1376 (.A(n_5_1269), .B1(n_5_1271), .B2(n_5_1318), .ZN(n_5_1233));
   OR2_X1 i_5_1377 (.A1(n_5_3168), .A2(n_55), .ZN(n_5_1234));
   NAND2_X1 i_5_1378 (.A1(n_5_3168), .A2(n_55), .ZN(n_5_1235));
   NAND2_X1 i_5_1393 (.A1(n_5_1234), .A2(n_5_1235), .ZN(n_5_1236));
   XNOR2_X1 i_5_1396 (.A(n_5_1233), .B(n_5_1236), .ZN(n_5_1951));
   NAND2_X1 i_5_1614 (.A1(n_5_1233), .A2(n_5_1234), .ZN(n_5_1237));
   NAND2_X1 i_5_1615 (.A1(n_5_1237), .A2(n_5_1235), .ZN(n_5_1238));
   XNOR2_X1 i_5_1616 (.A(n_5_3297), .B(n_73), .ZN(n_5_1239));
   XNOR2_X1 i_5_1617 (.A(n_5_1238), .B(n_5_1239), .ZN(n_5_1952));
   NAND2_X1 i_5_1618 (.A1(n_5_3297), .A2(n_73), .ZN(n_5_1240));
   XOR2_X1 i_5_1619 (.A(n_5_2017), .B(n_61), .Z(n_5_1241));
   NAND3_X1 i_5_1620 (.A1(n_5_1323), .A2(n_5_1324), .A3(n_5_1304), .ZN(n_5_1242));
   NAND2_X1 i_5_1621 (.A1(n_5_1242), .A2(n_5_1303), .ZN(n_5_1243));
   XNOR2_X1 i_5_1622 (.A(n_5_1241), .B(n_5_1243), .ZN(n_5_1954));
   NAND2_X1 i_5_1623 (.A1(n_5_2017), .A2(n_61), .ZN(n_5_1244));
   NAND2_X1 i_5_1624 (.A1(n_5_1221), .A2(n_5_1222), .ZN(n_5_1245));
   OAI21_X1 i_5_1625 (.A(n_5_1275), .B1(n_5_1274), .B2(n_5_1276), .ZN(n_5_1246));
   NAND2_X1 i_5_1626 (.A1(n_5_1246), .A2(n_5_1279), .ZN(n_5_2168));
   XNOR2_X1 i_5_1627 (.A(n_5_1227), .B(n_5_1219), .ZN(n_5_1247));
   BUF_X1 i_5_1628 (.A(n_5_1257), .Z(n_5_1248));
   BUF_X1 i_5_1629 (.A(n_5_1228), .Z(n_5_2169));
   BUF_X1 i_5_1630 (.A(n_5_1244), .Z(n_5_1249));
   BUF_X1 i_5_1631 (.A(n_5_1247), .Z(n_5_1250));
   NAND2_X1 i_5_1632 (.A1(n_5_464), .A2(n_53), .ZN(n_5_1251));
   NAND3_X1 i_5_1633 (.A1(n_5_1242), .A2(n_5_1245), .A3(n_5_1303), .ZN(n_5_1252));
   INV_X1 i_5_1634 (.A(n_5_1252), .ZN(n_5_1253));
   OAI211_X1 i_5_1635 (.A(n_5_1247), .B(n_5_1251), .C1(n_5_1253), .C2(n_5_1225), 
      .ZN(n_5_1254));
   INV_X1 i_5_1636 (.A(n_5_1250), .ZN(n_5_1255));
   NAND4_X1 i_5_1637 (.A1(n_5_1252), .A2(n_5_1255), .A3(n_5_1226), .A4(n_5_1249), 
      .ZN(n_5_1256));
   BUF_X1 i_5_1638 (.A(n_5_1251), .Z(n_5_1257));
   XNOR2_X1 i_5_1639 (.A(n_5_1784), .B(n_66), .ZN(n_5_2170));
   INV_X1 i_5_1640 (.A(n_5_1719), .ZN(n_5_1258));
   INV_X1 i_5_1641 (.A(n_58), .ZN(n_5_1259));
   NAND2_X1 i_5_1642 (.A1(n_5_3113), .A2(n_5_2866), .ZN(n_5_1260));
   OR2_X1 i_5_1643 (.A1(n_5_3113), .A2(n_5_2866), .ZN(n_5_1261));
   NAND2_X1 i_5_1644 (.A1(n_5_1287), .A2(n_5_1322), .ZN(n_5_1262));
   NAND2_X1 i_5_1645 (.A1(n_5_1302), .A2(n_5_2866), .ZN(n_5_1263));
   INV_X1 i_5_1397 (.A(n_5_1263), .ZN(n_5_1264));
   INV_X1 i_5_1647 (.A(n_5_2866), .ZN(n_5_1265));
   NAND2_X1 i_5_1408 (.A1(n_5_3028), .A2(n_5_1265), .ZN(n_5_1266));
   NOR2_X1 i_5_1410 (.A1(n_5_3028), .A2(n_5_1265), .ZN(n_5_1267));
   OAI21_X1 i_5_1415 (.A(n_5_1266), .B1(n_5_3113), .B2(n_5_1267), .ZN(n_5_1268));
   NOR2_X1 i_5_1416 (.A1(n_5_3137), .A2(n_60), .ZN(n_5_1269));
   INV_X1 i_5_1652 (.A(n_60), .ZN(n_5_1270));
   INV_X1 i_5_1438 (.A(n_5_1329), .ZN(n_5_1271));
   INV_X1 i_5_1654 (.A(n_5_1282), .ZN(n_5_1272));
   NAND2_X1 i_5_1655 (.A1(n_5_1240), .A2(n_5_1272), .ZN(n_5_1273));
   AND2_X1 i_5_1656 (.A1(n_5_1243), .A2(n_5_1244), .ZN(n_5_1274));
   XOR2_X1 i_5_1657 (.A(n_5_464), .B(n_53), .Z(n_5_1275));
   INV_X1 i_5_1658 (.A(n_5_1245), .ZN(n_5_1276));
   NAND2_X1 i_5_1659 (.A1(n_5_1243), .A2(n_5_1244), .ZN(n_5_1277));
   XNOR2_X1 i_5_1660 (.A(n_5_464), .B(n_53), .ZN(n_5_1278));
   NAND3_X1 i_5_1661 (.A1(n_5_1277), .A2(n_5_1278), .A3(n_5_1245), .ZN(n_5_1279));
   INV_X1 i_5_1662 (.A(n_66), .ZN(n_5_1280));
   NAND3_X1 i_5_1663 (.A1(n_5_1237), .A2(n_5_1235), .A3(n_5_1240), .ZN(n_5_1281));
   NAND2_X1 i_5_1664 (.A1(n_5_2936), .A2(n_5_1220), .ZN(n_5_1282));
   INV_X1 i_5_1665 (.A(n_5_1240), .ZN(n_5_1283));
   NAND2_X1 i_5_1666 (.A1(n_5_1237), .A2(n_5_1235), .ZN(n_5_1284));
   INV_X1 i_5_1667 (.A(n_58), .ZN(n_5_1285));
   NAND2_X1 i_5_1668 (.A1(n_5_1287), .A2(n_5_1322), .ZN(n_5_1286));
   NAND3_X1 i_5_1669 (.A1(n_5_1722), .A2(n_5_1327), .A3(n_5_1289), .ZN(n_5_1287));
   OR2_X1 i_5_1670 (.A1(n_5_2002), .A2(n_5_3329), .ZN(n_5_1288));
   NAND2_X1 i_5_1671 (.A1(n_5_2002), .A2(n_5_3329), .ZN(n_5_1289));
   XNOR2_X1 i_5_1672 (.A(n_5_2002), .B(n_5_3329), .ZN(n_5_1290));
   NAND2_X1 i_5_1673 (.A1(n_5_1254), .A2(n_5_1256), .ZN(n_5_1291));
   NOR2_X1 i_5_1674 (.A1(n_5_1248), .A2(n_5_1250), .ZN(n_5_1292));
   NOR2_X1 i_5_1675 (.A1(n_5_1291), .A2(n_5_1292), .ZN(n_5_1958));
   NAND2_X1 i_5_1676 (.A1(n_5_2963), .A2(n_5_3023), .ZN(n_5_1293));
   INV_X1 i_5_1677 (.A(n_5_1280), .ZN(n_5_1294));
   NOR2_X1 i_5_1678 (.A1(n_5_3185), .A2(n_5_1294), .ZN(n_5_1295));
   INV_X1 i_5_1679 (.A(n_5_1336), .ZN(n_5_1296));
   NAND2_X1 i_5_1680 (.A1(n_5_2963), .A2(n_5_1296), .ZN(n_5_1297));
   NAND3_X1 i_5_1681 (.A1(n_5_1334), .A2(n_5_1293), .A3(n_5_1297), .ZN(n_5_1298));
   NOR2_X1 i_5_1254 (.A1(n_5_1298), .A2(n_5_3093), .ZN(n_5_1959));
   INV_X1 i_5_1683 (.A(n_76), .ZN(n_5_1299));
   INV_X1 i_5_1684 (.A(n_5_3185), .ZN(n_5_1803));
   INV_X1 i_5_1685 (.A(n_5_1306), .ZN(n_5_1300));
   INV_X1 i_5_1686 (.A(n_5_2569), .ZN(n_5_1301));
   INV_X1 i_5_1687 (.A(n_5_2963), .ZN(n_5_1302));
   NAND2_X1 i_5_1688 (.A1(n_5_2948), .A2(n_5_1280), .ZN(n_5_3162));
   OR2_X1 i_5_1689 (.A1(n_5_2013), .A2(n_75), .ZN(n_5_1303));
   NAND2_X1 i_5_1690 (.A1(n_5_2013), .A2(n_75), .ZN(n_5_1304));
   INV_X1 i_5_1691 (.A(n_5_1331), .ZN(n_5_1305));
   NAND2_X1 i_5_1692 (.A1(n_5_1721), .A2(n_5_1289), .ZN(n_5_1306));
   NAND4_X1 i_5_1693 (.A1(n_5_3821), .A2(n_5_3106), .A3(n_5_1330), .A4(n_5_1268), 
      .ZN(n_5_1307));
   XNOR2_X1 i_5_1694 (.A(n_5_1321), .B(n_5_1307), .ZN(n_5_2174));
   INV_X1 i_5_1695 (.A(n_5_1280), .ZN(n_5_1308));
   NAND2_X1 i_5_1696 (.A1(n_5_1786), .A2(n_5_1308), .ZN(n_5_1309));
   INV_X1 i_5_1697 (.A(n_5_1786), .ZN(n_5_1310));
   OAI21_X1 i_5_1698 (.A(n_5_1309), .B1(n_5_2948), .B2(n_5_1310), .ZN(n_5_1311));
   XNOR2_X1 i_5_1699 (.A(n_5_1299), .B(n_5_1220), .ZN(n_5_1312));
   INV_X1 i_5_1700 (.A(n_5_1299), .ZN(n_5_1313));
   NAND2_X1 i_5_1701 (.A1(n_5_2936), .A2(n_5_1312), .ZN(n_5_1314));
   NAND2_X1 i_5_1702 (.A1(n_5_1312), .A2(n_5_1313), .ZN(n_5_1315));
   INV_X1 i_5_1703 (.A(n_5_2936), .ZN(n_5_1316));
   NAND2_X1 i_5_1704 (.A1(n_5_1316), .A2(n_5_1313), .ZN(n_5_1317));
   NAND2_X1 i_5_1439 (.A1(n_5_3137), .A2(n_60), .ZN(n_5_1318));
   INV_X1 i_5_1706 (.A(n_60), .ZN(n_5_1319));
   INV_X1 i_5_1707 (.A(n_5_1270), .ZN(n_5_1320));
   OAI22_X1 i_5_1708 (.A1(n_5_1755), .A2(n_5_1319), .B1(n_5_3137), .B2(n_5_1320), 
      .ZN(n_5_1321));
   OR2_X1 i_5_1709 (.A1(n_5_2012), .A2(n_5_2569), .ZN(n_5_1322));
   NAND3_X1 i_5_1710 (.A1(n_5_1325), .A2(n_5_1273), .A3(n_5_1281), .ZN(n_5_1323));
   NAND2_X1 i_5_1711 (.A1(n_5_1751), .A2(n_76), .ZN(n_5_1324));
   INV_X1 i_5_1712 (.A(n_5_1716), .ZN(n_5_3163));
   OR2_X1 i_5_1713 (.A1(n_5_1751), .A2(n_76), .ZN(n_5_1325));
   NAND2_X1 i_5_1714 (.A1(n_5_1288), .A2(n_5_1232), .ZN(n_5_1326));
   NAND2_X1 i_5_1715 (.A1(n_5_1326), .A2(n_5_1289), .ZN(n_5_2178));
   NAND2_X1 i_5_1716 (.A1(n_5_1288), .A2(n_5_1232), .ZN(n_5_1327));
   NAND2_X1 i_5_1457 (.A1(n_5_3112), .A2(n_5_1264), .ZN(n_5_1328));
   NAND4_X1 i_5_1467 (.A1(n_5_3821), .A2(n_5_3106), .A3(n_5_1328), .A4(n_5_1268), 
      .ZN(n_5_1329));
   NAND2_X1 i_5_1719 (.A1(n_5_3112), .A2(n_5_1264), .ZN(n_5_1330));
   INV_X1 i_5_1720 (.A(n_5_1262), .ZN(n_5_3164));
   NAND2_X1 i_5_1721 (.A1(n_5_1719), .A2(n_58), .ZN(n_5_1331));
   NAND3_X1 i_5_1722 (.A1(n_5_1785), .A2(n_5_3018), .A3(n_5_1786), .ZN(n_5_1332));
   AOI22_X1 i_5_1723 (.A1(n_5_1784), .A2(n_66), .B1(n_5_1719), .B2(n_58), 
      .ZN(n_5_1333));
   NAND3_X1 i_5_1724 (.A1(n_5_3026), .A2(n_5_1332), .A3(n_5_1333), .ZN(n_5_1334));
   INV_X1 i_5_1725 (.A(n_5_1784), .ZN(n_5_1335));
   NAND2_X1 i_5_1726 (.A1(n_5_1335), .A2(n_5_1295), .ZN(n_5_1336));
   NAND2_X1 i_5_1727 (.A1(n_5_2948), .A2(n_5_1280), .ZN(n_5_1964));
   NAND2_X1 i_5_1728 (.A1(n_5_1335), .A2(n_5_1280), .ZN(n_5_1337));
   NAND2_X1 i_5_1729 (.A1(n_5_2948), .A2(n_5_1280), .ZN(n_5_1338));
   INV_X1 i_5_1730 (.A(m[14]), .ZN(n_5_1339));
   INV_X1 i_5_1731 (.A(m[15]), .ZN(n_5_1340));
   NAND2_X1 i_5_1732 (.A1(n_5_1429), .A2(m[0]), .ZN(n_5_1341));
   INV_X1 i_5_1733 (.A(m[1]), .ZN(n_5_1342));
   INV_X1 i_5_1734 (.A(m[2]), .ZN(n_5_1966));
   INV_X1 i_5_1735 (.A(m[3]), .ZN(n_5_1967));
   INV_X1 i_5_1736 (.A(m[4]), .ZN(n_5_2179));
   INV_X1 i_5_1737 (.A(m[5]), .ZN(n_5_2180));
   INV_X1 i_5_1738 (.A(m[6]), .ZN(n_5_2181));
   INV_X1 i_5_1739 (.A(m[7]), .ZN(n_5_1343));
   INV_X1 i_5_1740 (.A(n_5_3137), .ZN(n_5_1969));
   INV_X1 i_5_1741 (.A(m[8]), .ZN(n_5_1970));
   NAND2_X1 i_5_1742 (.A1(n_5_3137), .A2(m[8]), .ZN(n_5_3165));
   INV_X1 i_5_1743 (.A(n_5_3168), .ZN(n_5_3166));
   INV_X1 i_5_1744 (.A(m[9]), .ZN(n_5_3167));
   INV_X1 i_5_1745 (.A(m[10]), .ZN(n_5_1344));
   NAND2_X1 i_5_1746 (.A1(n_5_2970), .A2(n_5_1344), .ZN(n_5_1345));
   INV_X1 i_5_1747 (.A(m[11]), .ZN(n_5_1971));
   INV_X1 i_5_1748 (.A(m[12]), .ZN(n_5_1346));
   NAND2_X1 i_5_1749 (.A1(n_5_1732), .A2(n_5_1346), .ZN(n_5_1347));
   INV_X1 i_5_1750 (.A(n_5_2017), .ZN(n_5_1348));
   INV_X1 i_5_1751 (.A(m[13]), .ZN(n_5_1349));
   NAND2_X1 i_5_1752 (.A1(n_5_1348), .A2(n_5_1349), .ZN(n_5_1350));
   NAND2_X1 i_5_1753 (.A1(n_5_464), .A2(m[14]), .ZN(n_5_1351));
   INV_X1 i_5_1754 (.A(n_5_464), .ZN(n_5_1352));
   NAND2_X1 i_5_1755 (.A1(n_5_1352), .A2(n_5_1339), .ZN(n_5_1353));
   OAI21_X1 i_5_1756 (.A(n_5_2999), .B1(n_5_1341), .B2(n_5_1356), .ZN(n_5_1354));
   NAND3_X1 i_5_1757 (.A1(n_5_1414), .A2(n_5_1341), .A3(n_5_2999), .ZN(n_5_1355));
   INV_X1 i_5_1758 (.A(n_5_1410), .ZN(n_5_1356));
   NAND2_X1 i_5_1759 (.A1(n_5_1414), .A2(n_5_1356), .ZN(n_5_1357));
   NAND3_X1 i_5_1760 (.A1(n_5_1355), .A2(n_5_1357), .A3(n_5_2997), .ZN(n_5_1358));
   AOI21_X1 i_5_1761 (.A(n_5_3238), .B1(n_5_1416), .B2(n_5_1527), .ZN(n_5_2182));
   INV_X1 i_5_1255 (.A(n_5_1542), .ZN(n_5_1359));
   NAND3_X1 i_5_1256 (.A1(n_5_3025), .A2(n_5_1530), .A3(n_5_1359), .ZN(n_5_1360));
   INV_X1 i_5_1764 (.A(n_5_3454), .ZN(n_5_1361));
   OAI21_X1 i_5_1257 (.A(n_5_3354), .B1(n_5_1361), .B2(n_5_1527), .ZN(n_5_1362));
   NAND2_X1 i_5_1262 (.A1(n_5_3025), .A2(n_5_1362), .ZN(n_5_1363));
   NAND3_X1 i_5_1263 (.A1(n_5_1360), .A2(n_5_1363), .A3(n_5_1528), .ZN(n_5_1364));
   INV_X1 i_5_1768 (.A(n_5_1386), .ZN(n_5_1365));
   NAND2_X1 i_5_1769 (.A1(n_5_2937), .A2(n_5_3165), .ZN(n_5_1366));
   NAND2_X1 i_5_1770 (.A1(n_5_1560), .A2(n_5_1345), .ZN(n_5_1367));
   NAND2_X1 i_5_1771 (.A1(n_5_3532), .A2(n_5_1529), .ZN(n_5_1368));
   INV_X1 i_5_1772 (.A(n_5_1345), .ZN(n_5_1369));
   AOI21_X1 i_5_1773 (.A(n_5_3473), .B1(n_5_1365), .B2(n_5_1416), .ZN(n_5_1370));
   INV_X1 i_5_1774 (.A(n_5_1733), .ZN(n_5_1371));
   NAND3_X1 i_5_1775 (.A1(n_5_1399), .A2(n_5_1779), .A3(n_5_1733), .ZN(n_5_1372));
   NAND3_X1 i_5_1342 (.A1(n_5_1372), .A2(n_5_1782), .A3(n_5_1350), .ZN(n_5_461));
   NAND2_X1 i_5_1778 (.A1(n_5_1779), .A2(n_5_1733), .ZN(n_5_1375));
   INV_X1 i_5_1779 (.A(n_5_1375), .ZN(n_5_1376));
   NAND2_X1 i_5_1780 (.A1(n_5_1350), .A2(n_5_1347), .ZN(n_5_1377));
   NAND3_X1 i_5_1781 (.A1(n_5_1377), .A2(n_5_1353), .A3(n_5_1779), .ZN(n_5_1378));
   NAND3_X1 i_5_1782 (.A1(n_5_1396), .A2(n_5_1378), .A3(n_5_1351), .ZN(n_5_1972));
   XNOR2_X1 i_5_1783 (.A(n_5_2006), .B(m[1]), .ZN(n_5_1379));
   XNOR2_X1 i_5_1784 (.A(n_5_1409), .B(n_5_1379), .ZN(n_5_1973));
   XNOR2_X1 i_5_1785 (.A(n_5_2002), .B(m[2]), .ZN(n_5_1380));
   XNOR2_X1 i_5_1786 (.A(n_5_1380), .B(n_5_1354), .ZN(n_5_1974));
   XNOR2_X1 i_5_1787 (.A(n_5_1531), .B(n_5_1783), .ZN(n_5_3387));
   XNOR2_X1 i_5_1788 (.A(n_5_2017), .B(m[13]), .ZN(n_5_1381));
   XNOR2_X1 i_5_1789 (.A(n_5_1420), .B(n_5_1381), .ZN(n_5_1977));
   XNOR2_X1 i_5_1792 (.A(n_5_1340), .B(m[14]), .ZN(n_5_1979));
   NAND2_X1 i_5_1793 (.A1(n_5_1765), .A2(n_5_3025), .ZN(n_5_1383));
   INV_X1 i_5_1794 (.A(n_5_3165), .ZN(n_5_1384));
   INV_X1 i_5_1795 (.A(m[10]), .ZN(n_5_1385));
   AND2_X1 i_5_1796 (.A1(n_5_1421), .A2(n_5_1573), .ZN(n_5_2185));
   BUF_X1 i_5_1797 (.A(n_5_1392), .Z(n_5_1386));
   INV_X1 i_5_1798 (.A(m[3]), .ZN(n_5_1387));
   XNOR2_X1 i_5_1799 (.A(n_5_1358), .B(n_5_1724), .ZN(n_5_1980));
   INV_X1 i_5_1800 (.A(n_5_2938), .ZN(n_5_1388));
   INV_X1 i_5_1801 (.A(n_5_2939), .ZN(n_5_1389));
   INV_X1 i_5_1802 (.A(n_5_2940), .ZN(n_5_1390));
   NAND2_X1 i_5_1803 (.A1(n_5_2185), .A2(n_5_1400), .ZN(n_5_2186));
   NAND2_X1 i_5_1804 (.A1(n_5_1369), .A2(n_5_1424), .ZN(n_5_1982));
   OAI211_X1 i_5_1776 (.A(n_5_1424), .B(n_5_3535), .C1(n_5_1370), .C2(n_5_1368), 
      .ZN(n_5_1983));
   AOI22_X1 i_5_1777 (.A1(n_5_1550), .A2(n_5_1383), .B1(m[7]), .B2(n_5_3113), 
      .ZN(n_5_1391));
   NAND2_X1 i_5_1807 (.A1(n_5_1417), .A2(n_5_1550), .ZN(n_5_1392));
   NAND2_X1 i_5_1808 (.A1(n_5_3113), .A2(m[7]), .ZN(n_5_2187));
   INV_X1 i_5_1809 (.A(n_5_1532), .ZN(n_5_1393));
   AOI21_X1 i_5_1810 (.A(n_5_1383), .B1(n_5_1417), .B2(n_5_1393), .ZN(n_5_2188));
   INV_X1 i_5_1811 (.A(m[7]), .ZN(n_5_1394));
   XNOR2_X1 i_5_1266 (.A(n_5_3113), .B(n_5_1394), .ZN(n_5_1395));
   XNOR2_X1 i_5_1273 (.A(n_5_1364), .B(n_5_1395), .ZN(n_5_1984));
   NAND4_X1 i_5_1814 (.A1(n_5_1376), .A2(n_5_1399), .A3(n_5_1353), .A4(n_5_1350), 
      .ZN(n_5_1396));
   NAND2_X1 i_5_1815 (.A1(n_5_3010), .A2(n_5_3009), .ZN(n_5_1397));
   NAND2_X1 i_5_1816 (.A1(n_5_3011), .A2(n_5_3009), .ZN(n_5_1398));
   NAND2_X1 i_5_1817 (.A1(n_5_1397), .A2(n_5_1398), .ZN(n_5_1399));
   OAI22_X1 i_5_1818 (.A1(n_5_1401), .A2(m[10]), .B1(n_5_3297), .B2(n_5_1385), 
      .ZN(n_5_1400));
   INV_X1 i_5_1819 (.A(n_5_3297), .ZN(n_5_1401));
   INV_X1 i_5_1820 (.A(n_5_1385), .ZN(n_5_1402));
   XNOR2_X1 i_5_1821 (.A(n_5_3532), .B(n_5_1402), .ZN(n_5_1403));
   INV_X1 i_5_1822 (.A(n_5_3297), .ZN(n_5_1404));
   NAND2_X1 i_5_1823 (.A1(n_5_1403), .A2(n_5_1404), .ZN(n_5_1405));
   INV_X1 i_5_1824 (.A(m[10]), .ZN(n_5_1406));
   XNOR2_X1 i_5_1825 (.A(n_5_3532), .B(n_5_1406), .ZN(n_5_1407));
   NAND2_X1 i_5_1826 (.A1(n_5_1407), .A2(n_5_3297), .ZN(n_5_1408));
   NAND2_X1 i_5_1827 (.A1(n_5_1405), .A2(n_5_1408), .ZN(n_5_2189));
   INV_X1 i_5_1828 (.A(n_5_1341), .ZN(n_5_1409));
   NAND2_X1 i_5_1829 (.A1(n_5_1565), .A2(n_5_1342), .ZN(n_5_1410));
   NAND2_X1 i_5_1830 (.A1(n_5_1565), .A2(n_5_1342), .ZN(n_5_1411));
   INV_X1 i_5_1831 (.A(n_5_1411), .ZN(n_5_1412));
   INV_X1 i_5_1832 (.A(m[5]), .ZN(n_5_1413));
   XNOR2_X1 i_5_1833 (.A(n_5_1784), .B(n_5_1413), .ZN(n_5_2190));
   NAND2_X1 i_5_1834 (.A1(n_5_2002), .A2(m[2]), .ZN(n_5_1414));
   NAND2_X1 i_5_1835 (.A1(n_5_2002), .A2(m[2]), .ZN(n_5_1986));
   OAI21_X1 i_5_1836 (.A(n_5_1388), .B1(n_5_1389), .B2(n_5_1390), .ZN(n_5_1415));
   XNOR2_X1 i_5_1837 (.A(n_5_1415), .B(n_5_1718), .ZN(n_5_1987));
   OAI21_X1 i_5_1838 (.A(n_5_1388), .B1(n_5_1389), .B2(n_5_1390), .ZN(n_5_1416));
   AOI21_X1 i_5_1839 (.A(n_5_3369), .B1(n_5_3314), .B2(n_5_2181), .ZN(n_5_1417));
   NAND2_X1 i_5_1840 (.A1(n_5_3190), .A2(n_5_1347), .ZN(n_5_1418));
   INV_X1 i_5_1841 (.A(n_5_1371), .ZN(n_5_1419));
   NAND2_X1 i_5_1842 (.A1(n_5_1418), .A2(n_5_1419), .ZN(n_5_1420));
   OAI21_X1 i_5_1843 (.A(n_5_2974), .B1(n_5_1384), .B2(n_5_2025), .ZN(n_5_1421));
   INV_X1 i_5_1844 (.A(m[9]), .ZN(n_5_1988));
   NOR2_X1 i_5_1845 (.A1(n_5_2025), .A2(n_5_1384), .ZN(n_5_1422));
   NAND2_X1 i_5_1479 (.A1(n_5_2973), .A2(n_5_1422), .ZN(n_5_1423));
   OAI21_X1 i_5_1573 (.A(n_5_1423), .B1(n_5_2982), .B2(n_5_1422), .ZN(n_5_1989));
   NAND2_X1 i_5_1848 (.A1(n_5_3297), .A2(m[10]), .ZN(n_5_1424));
   NAND2_X1 i_5_1849 (.A1(n_5_1462), .A2(n_5_3170), .ZN(n_5_1425));
   NAND2_X1 i_5_1850 (.A1(n_5_1812), .A2(n_5_1453), .ZN(n_5_1426));
   INV_X1 i_5_1851 (.A(n_5_1426), .ZN(n_5_1427));
   AOI21_X1 i_5_1852 (.A(n_5_1427), .B1(n_5_1587), .B2(n_5_1452), .ZN(n_5_1428));
   NAND2_X1 i_5_1853 (.A1(n_5_1425), .A2(n_5_1428), .ZN(n_5_1429));
   NAND2_X1 i_5_1854 (.A1(n_5_1465), .A2(n_5_3170), .ZN(n_5_1430));
   NAND2_X1 i_5_1855 (.A1(n_5_3822), .A2(n_5_1453), .ZN(n_5_1431));
   NAND2_X1 i_5_1856 (.A1(n_5_1592), .A2(n_5_1452), .ZN(n_5_1432));
   NAND2_X1 i_5_1857 (.A1(n_5_1467), .A2(n_5_3170), .ZN(n_5_1433));
   NAND2_X1 i_5_1858 (.A1(n_5_2918), .A2(n_5_1453), .ZN(n_5_1434));
   NAND2_X1 i_5_1859 (.A1(n_5_3348), .A2(n_5_1453), .ZN(n_5_1435));
   NAND2_X1 i_5_1860 (.A1(n_5_3554), .A2(n_5_1453), .ZN(n_5_1436));
   NAND2_X1 i_5_1861 (.A1(n_5_1499), .A2(n_5_3170), .ZN(n_5_1437));
   NAND2_X1 i_5_1862 (.A1(n_5_1602), .A2(n_5_1452), .ZN(n_5_1438));
   NAND2_X1 i_5_1863 (.A1(n_5_3412), .A2(n_5_1453), .ZN(n_5_1439));
   NAND2_X1 i_5_1579 (.A1(n_5_3733), .A2(n_5_1453), .ZN(n_5_2191));
   NAND2_X1 i_5_1865 (.A1(n_5_1816), .A2(n_5_1453), .ZN(n_5_2192));
   NAND2_X1 i_5_1866 (.A1(n_5_3094), .A2(n_5_1453), .ZN(n_5_1440));
   NAND2_X1 i_5_1867 (.A1(n_5_3107), .A2(n_5_1453), .ZN(n_5_1441));
   NAND3_X1 i_5_1580 (.A1(n_5_1789), .A2(n_5_1726), .A3(n_5_1441), .ZN(n_5_3168));
   NAND2_X1 i_5_1869 (.A1(n_5_4462), .A2(n_5_1453), .ZN(n_5_1442));
   NAND2_X1 i_5_1870 (.A1(n_5_1821), .A2(n_5_1453), .ZN(n_5_1443));
   INV_X1 i_5_1871 (.A(n_5_1443), .ZN(n_5_1444));
   AOI21_X1 i_5_1872 (.A(n_5_1444), .B1(n_5_1603), .B2(n_5_1452), .ZN(n_5_1445));
   NAND2_X1 i_5_1873 (.A1(n_5_1470), .A2(n_5_3170), .ZN(n_5_1446));
   NAND2_X1 i_5_1874 (.A1(n_5_3191), .A2(n_5_1453), .ZN(n_5_1447));
   INV_X1 i_5_1875 (.A(n_5_1447), .ZN(n_5_1448));
   AOI21_X1 i_5_1876 (.A(n_5_1448), .B1(n_5_1664), .B2(n_5_1452), .ZN(n_5_1449));
   INV_X1 i_5_1877 (.A(r[2]), .ZN(n_5_1450));
   NAND2_X1 i_5_1878 (.A1(r[3]), .A2(n_5_1450), .ZN(n_5_1451));
   INV_X1 i_5_1879 (.A(n_5_1451), .ZN(n_5_1452));
   NOR2_X1 i_5_1880 (.A1(r[3]), .A2(n_5_1450), .ZN(n_5_3170));
   XNOR2_X1 i_5_1881 (.A(r[3]), .B(r[2]), .ZN(n_5_1453));
   NAND2_X1 i_5_1882 (.A1(n_5_3246), .A2(n_5_1453), .ZN(n_5_3171));
   NAND2_X1 i_5_1883 (.A1(n_5_1622), .A2(n_5_1452), .ZN(n_5_1454));
   INV_X1 i_5_1884 (.A(n_5_1442), .ZN(n_5_2196));
   NAND2_X1 i_5_1885 (.A1(n_5_1469), .A2(n_5_3170), .ZN(n_5_1455));
   NAND2_X1 i_5_1886 (.A1(n_5_1621), .A2(n_5_1452), .ZN(n_5_1456));
   NAND2_X1 i_5_1887 (.A1(n_5_1775), .A2(n_5_3170), .ZN(n_5_1457));
   NAND2_X1 i_5_1274 (.A1(n_5_1468), .A2(n_5_3170), .ZN(n_5_2197));
   NAND2_X1 i_5_1275 (.A1(n_5_1666), .A2(n_5_1452), .ZN(n_5_2198));
   NAND2_X1 i_5_1890 (.A1(n_5_3374), .A2(n_5_3525), .ZN(n_5_2199));
   NAND2_X1 i_5_1891 (.A1(n_5_3449), .A2(n_5_4218), .ZN(n_5_3172));
   INV_X1 i_5_1892 (.A(n_5_1458), .ZN(n_5_4065));
   XNOR2_X1 i_5_1893 (.A(n_5_1459), .B(m[14]), .ZN(n_5_1458));
   INV_X1 i_5_1894 (.A(m[15]), .ZN(n_5_1459));
   NAND2_X1 i_5_1895 (.A1(n_5_3246), .A2(m[14]), .ZN(n_5_1460));
   INV_X1 i_5_1896 (.A(m[9]), .ZN(n_5_1461));
   INV_X1 i_5_1897 (.A(n_5_3191), .ZN(n_5_3173));
   INV_X1 i_5_1898 (.A(m[13]), .ZN(n_5_3174));
   INV_X1 i_5_1899 (.A(n_5_2204), .ZN(n_5_2202));
   XOR2_X1 i_5_1900 (.A(n_5_1494), .B(n_5_1463), .Z(n_5_1462));
   OR2_X1 i_5_1901 (.A1(n_5_1464), .A2(n_5_1493), .ZN(n_5_1463));
   INV_X1 i_5_1902 (.A(n_5_1511), .ZN(n_5_1464));
   XNOR2_X1 i_5_1903 (.A(n_5_1466), .B(n_5_1512), .ZN(n_5_1465));
   NAND2_X1 i_5_1904 (.A1(n_5_3824), .A2(n_5_1473), .ZN(n_5_1466));
   XOR2_X1 i_5_1905 (.A(n_5_1503), .B(n_5_1492), .Z(n_5_1467));
   XOR2_X1 i_5_1291 (.A(n_5_1571), .B(n_5_1501), .Z(n_5_1468));
   OAI21_X1 i_5_1907 (.A(n_5_1540), .B1(n_5_3477), .B2(n_5_1533), .ZN(n_5_2203));
   XOR2_X1 i_5_1908 (.A(n_5_3485), .B(n_5_1557), .Z(n_5_1469));
   XOR2_X1 i_5_1909 (.A(n_5_3529), .B(n_5_2206), .Z(n_5_1470));
   NAND2_X1 i_5_1910 (.A1(n_5_4085), .A2(n_5_1460), .ZN(n_5_2204));
   NAND2_X1 i_5_1911 (.A1(n_5_1471), .A2(n_5_1555), .ZN(n_5_2206));
   NAND2_X1 i_5_1912 (.A1(n_5_3485), .A2(n_5_1556), .ZN(n_5_1471));
   INV_X1 i_5_1913 (.A(n_5_3102), .ZN(n_5_3175));
   INV_X1 i_5_1914 (.A(n_5_1473), .ZN(n_5_1472));
   NAND2_X1 i_5_1915 (.A1(n_5_3822), .A2(m[2]), .ZN(n_5_1473));
   NAND2_X1 i_5_1916 (.A1(n_5_4462), .A2(m[11]), .ZN(n_5_3176));
   NOR2_X1 i_5_1917 (.A1(n_5_3412), .A2(m[6]), .ZN(n_5_1474));
   INV_X1 i_5_1918 (.A(m[6]), .ZN(n_5_1475));
   OR2_X1 i_5_1919 (.A1(n_5_3733), .A2(m[7]), .ZN(n_5_1476));
   AOI21_X1 i_5_1612 (.A(n_5_1474), .B1(n_5_1514), .B2(n_5_1516), .ZN(n_5_2000));
   INV_X1 i_5_1921 (.A(n_5_3733), .ZN(n_5_1477));
   INV_X1 i_5_1922 (.A(m[7]), .ZN(n_5_1478));
   OR2_X1 i_5_1923 (.A1(n_5_3348), .A2(m[4]), .ZN(n_5_1479));
   NAND2_X1 i_5_1646 (.A1(n_5_1476), .A2(n_5_1480), .ZN(n_5_2001));
   NAND2_X1 i_5_1925 (.A1(n_5_3733), .A2(m[7]), .ZN(n_5_1480));
   NAND2_X1 i_5_1926 (.A1(n_5_1571), .A2(n_5_1500), .ZN(n_5_2207));
   NAND2_X1 i_5_1927 (.A1(n_5_3094), .A2(m[9]), .ZN(n_5_1481));
   INV_X1 i_5_1928 (.A(m[8]), .ZN(n_5_1482));
   XNOR2_X1 i_5_1929 (.A(n_5_1461), .B(n_5_1482), .ZN(n_5_1483));
   MUX2_X1 i_5_1930 (.A(n_5_1461), .B(n_5_1483), .S(n_5_1816), .Z(n_5_2208));
   XNOR2_X1 i_5_1931 (.A(n_5_1482), .B(m[9]), .ZN(n_5_1484));
   MUX2_X1 i_5_1932 (.A(m[9]), .B(n_5_1484), .S(n_5_1816), .Z(n_5_2209));
   INV_X1 i_5_1933 (.A(n_5_1816), .ZN(n_5_1485));
   NAND2_X1 i_5_1934 (.A1(n_5_1485), .A2(n_5_1482), .ZN(n_5_1486));
   NAND4_X1 i_5_1935 (.A1(n_5_1486), .A2(n_5_1566), .A3(n_5_1567), .A4(n_5_1568), 
      .ZN(n_5_1487));
   INV_X1 i_5_1936 (.A(n_5_1487), .ZN(n_5_1488));
   INV_X1 i_5_1937 (.A(n_5_1461), .ZN(n_5_1489));
   INV_X1 i_5_1938 (.A(m[9]), .ZN(n_5_1490));
   MUX2_X1 i_5_1939 (.A(n_5_1489), .B(n_5_1490), .S(n_5_3094), .Z(n_5_1491));
   NAND2_X1 i_5_1940 (.A1(n_5_2917), .A2(n_5_2915), .ZN(n_5_1492));
   NOR2_X1 i_5_1941 (.A1(n_5_1812), .A2(m[1]), .ZN(n_5_1493));
   NAND2_X1 i_5_1942 (.A1(n_5_1811), .A2(m[0]), .ZN(n_5_1494));
   NAND3_X1 i_5_1943 (.A1(n_5_1812), .A2(n_5_1811), .A3(m[0]), .ZN(n_5_1495));
   NAND2_X1 i_5_1944 (.A1(m[0]), .A2(m[1]), .ZN(n_5_1496));
   INV_X1 i_5_1945 (.A(n_5_1496), .ZN(n_5_1497));
   NAND2_X1 i_5_1946 (.A1(n_5_1811), .A2(n_5_1497), .ZN(n_5_1498));
   XNOR2_X1 i_5_1947 (.A(n_5_1507), .B(n_5_1773), .ZN(n_5_1499));
   OR2_X1 i_5_1948 (.A1(n_5_1816), .A2(m[8]), .ZN(n_5_2210));
   NAND2_X1 i_5_1949 (.A1(n_5_1816), .A2(m[8]), .ZN(n_5_1500));
   XNOR2_X1 i_5_1292 (.A(n_5_1816), .B(m[8]), .ZN(n_5_1501));
   OAI21_X1 i_5_1951 (.A(n_5_3824), .B1(n_5_1513), .B2(n_5_1472), .ZN(n_5_1502));
   NAND2_X1 i_5_1952 (.A1(n_5_2915), .A2(n_5_1502), .ZN(n_5_1804));
   OAI21_X1 i_5_1953 (.A(n_5_3824), .B1(n_5_1513), .B2(n_5_1472), .ZN(n_5_1503));
   INV_X1 i_5_1954 (.A(n_5_3412), .ZN(n_5_1504));
   INV_X1 i_5_1955 (.A(m[6]), .ZN(n_5_1505));
   INV_X1 i_5_1956 (.A(n_5_1475), .ZN(n_5_1506));
   OAI22_X1 i_5_1957 (.A1(n_5_1504), .A2(n_5_1505), .B1(n_5_3412), .B2(n_5_1506), 
      .ZN(n_5_1507));
   INV_X1 i_5_1958 (.A(n_5_3183), .ZN(n_5_1508));
   INV_X1 i_5_1959 (.A(n_5_1762), .ZN(n_5_1509));
   NAND2_X1 i_5_1960 (.A1(n_5_1508), .A2(n_5_1509), .ZN(n_5_3177));
   NAND2_X1 i_5_1961 (.A1(n_5_1812), .A2(m[1]), .ZN(n_5_1510));
   NAND2_X1 i_5_1962 (.A1(n_5_1812), .A2(m[1]), .ZN(n_5_1511));
   AOI21_X1 i_5_1963 (.A(n_5_1493), .B1(n_5_1510), .B2(n_5_1494), .ZN(n_5_1512));
   NAND3_X1 i_5_1964 (.A1(n_5_1495), .A2(n_5_1510), .A3(n_5_1498), .ZN(n_5_1513));
   INV_X1 i_5_1965 (.A(n_5_1774), .ZN(n_5_1514));
   NAND2_X1 i_5_1966 (.A1(n_5_3733), .A2(m[7]), .ZN(n_5_1515));
   NAND2_X1 i_5_1967 (.A1(n_5_3412), .A2(m[6]), .ZN(n_5_1516));
   NAND2_X1 i_5_1968 (.A1(n_5_3412), .A2(m[6]), .ZN(n_5_1517));
   NAND3_X1 i_5_1969 (.A1(n_5_1517), .A2(n_5_1772), .A3(n_5_3551), .ZN(n_5_1518));
   NAND2_X1 i_5_1970 (.A1(n_5_1517), .A2(n_5_3550), .ZN(n_5_1519));
   NAND2_X1 i_5_1971 (.A1(n_5_1518), .A2(n_5_1519), .ZN(n_5_1520));
   NAND2_X1 i_5_1972 (.A1(n_5_3733), .A2(m[7]), .ZN(n_5_1521));
   NAND3_X1 i_5_1973 (.A1(n_5_1432), .A2(n_5_1433), .A3(n_5_1434), .ZN(n_5_2002));
   NAND3_X1 i_5_1974 (.A1(n_5_1433), .A2(n_5_1432), .A3(n_5_1434), .ZN(n_5_2003));
   NAND2_X1 i_5_1975 (.A1(n_5_3168), .A2(m[9]), .ZN(n_5_1522));
   INV_X1 i_5_1976 (.A(n_5_1522), .ZN(n_5_1523));
   NAND2_X1 i_5_1977 (.A1(n_5_1804), .A2(n_5_2916), .ZN(n_5_1524));
   NAND2_X1 i_5_1978 (.A1(n_5_1524), .A2(n_5_3344), .ZN(n_5_1525));
   NAND2_X1 i_5_1979 (.A1(n_5_2947), .A2(m[5]), .ZN(n_5_1526));
   NAND2_X1 i_5_1980 (.A1(n_5_3362), .A2(n_5_2179), .ZN(n_5_1527));
   NAND2_X1 i_5_1295 (.A1(n_5_3314), .A2(n_5_2181), .ZN(n_5_1528));
   NAND2_X1 i_5_1982 (.A1(n_5_1969), .A2(n_5_1970), .ZN(n_5_1529));
   BUF_X1 i_5_1296 (.A(n_5_2945), .Z(n_5_1530));
   AOI21_X1 i_5_1984 (.A(n_5_3021), .B1(n_5_1545), .B2(n_5_2945), .ZN(n_5_1531));
   AOI21_X1 i_5_1985 (.A(n_5_2938), .B1(n_5_2939), .B2(n_5_2940), .ZN(n_5_1532));
   NOR2_X1 i_5_1986 (.A1(n_5_4462), .A2(m[11]), .ZN(n_5_1533));
   NAND2_X1 i_5_1987 (.A1(n_5_3175), .A2(n_5_1762), .ZN(n_5_1534));
   INV_X1 i_5_1988 (.A(n_5_4462), .ZN(n_5_1535));
   INV_X1 i_5_1989 (.A(m[11]), .ZN(n_5_1536));
   NAND2_X1 i_5_1990 (.A1(n_5_1535), .A2(n_5_1536), .ZN(n_5_1537));
   NAND2_X1 i_5_1991 (.A1(n_5_3176), .A2(n_5_1537), .ZN(n_5_1538));
   INV_X1 i_5_1992 (.A(n_5_3183), .ZN(n_5_1539));
   NAND3_X1 i_5_1993 (.A1(n_5_1534), .A2(n_5_1538), .A3(n_5_1539), .ZN(n_5_1540));
   NAND2_X1 i_5_1994 (.A1(n_5_1719), .A2(m[4]), .ZN(n_5_1541));
   NAND3_X1 i_5_1995 (.A1(n_5_3454), .A2(n_5_1527), .A3(n_5_3239), .ZN(n_5_1542));
   INV_X1 i_5_1996 (.A(n_5_3358), .ZN(n_5_1543));
   NAND2_X1 i_5_1997 (.A1(n_5_1541), .A2(n_5_3454), .ZN(n_5_1544));
   NOR2_X1 i_5_1998 (.A1(n_5_1543), .A2(n_5_1544), .ZN(n_5_1545));
   NAND2_X1 i_5_1999 (.A1(n_5_3532), .A2(n_5_1529), .ZN(n_5_1546));
   INV_X1 i_5_2000 (.A(n_5_1546), .ZN(n_5_1547));
   NAND2_X1 i_5_2001 (.A1(n_5_2998), .A2(n_5_1966), .ZN(n_5_1548));
   NOR2_X1 i_5_2002 (.A1(n_5_1412), .A2(n_5_1341), .ZN(n_5_1549));
   NAND2_X1 i_5_2003 (.A1(n_5_1548), .A2(n_5_1549), .ZN(n_5_2004));
   NAND2_X1 i_5_2004 (.A1(n_5_1563), .A2(n_5_1343), .ZN(n_5_1550));
   NAND2_X1 i_5_2005 (.A1(n_5_1563), .A2(n_5_1343), .ZN(n_5_1551));
   INV_X1 i_5_2006 (.A(n_5_1551), .ZN(n_5_2211));
   INV_X1 i_5_2007 (.A(n_5_1487), .ZN(n_5_1552));
   NAND2_X1 i_5_2008 (.A1(n_5_1552), .A2(n_5_3170), .ZN(n_5_1553));
   OAI21_X1 i_5_2009 (.A(n_5_1440), .B1(n_5_1553), .B2(n_5_1491), .ZN(n_5_2212));
   INV_X1 i_5_2010 (.A(n_5_3170), .ZN(n_5_1554));
   NOR2_X1 i_5_2011 (.A1(n_5_1488), .A2(n_5_1554), .ZN(n_5_2213));
   OR2_X1 i_5_2012 (.A1(n_5_1821), .A2(m[12]), .ZN(n_5_1555));
   NAND2_X1 i_5_2013 (.A1(n_5_1821), .A2(m[12]), .ZN(n_5_1556));
   XNOR2_X1 i_5_2014 (.A(n_5_1821), .B(m[12]), .ZN(n_5_1557));
   NAND2_X1 i_5_2015 (.A1(n_5_1366), .A2(n_5_1547), .ZN(n_5_1558));
   AOI21_X1 i_5_2016 (.A(n_5_1523), .B1(n_5_3297), .B2(m[10]), .ZN(n_5_1559));
   NAND2_X1 i_5_2017 (.A1(n_5_1558), .A2(n_5_1559), .ZN(n_5_1560));
   NAND3_X1 i_5_2018 (.A1(n_5_1767), .A2(n_5_1766), .A3(n_5_3171), .ZN(n_5_1561));
   NAND3_X1 i_5_1790 (.A1(n_5_2197), .A2(n_5_2198), .A3(n_5_2192), .ZN(n_5_1562));
   INV_X1 i_5_1791 (.A(n_5_1562), .ZN(n_5_1563));
   NAND3_X1 i_5_2021 (.A1(n_5_3917), .A2(n_5_1430), .A3(n_5_1431), .ZN(n_5_2006));
   NAND3_X1 i_5_2022 (.A1(n_5_3917), .A2(n_5_1430), .A3(n_5_1431), .ZN(n_5_1564));
   INV_X1 i_5_2023 (.A(n_5_1564), .ZN(n_5_1565));
   NAND2_X1 i_5_2024 (.A1(n_5_1520), .A2(n_5_1521), .ZN(n_5_1566));
   NAND2_X1 i_5_2025 (.A1(n_5_1515), .A2(n_5_1474), .ZN(n_5_1567));
   NAND2_X1 i_5_2026 (.A1(n_5_1477), .A2(n_5_1478), .ZN(n_5_1568));
   NAND2_X1 i_5_2027 (.A1(n_5_1520), .A2(n_5_1521), .ZN(n_5_1569));
   AOI22_X1 i_5_2028 (.A1(n_5_1515), .A2(n_5_1474), .B1(n_5_1477), .B2(n_5_1478), 
      .ZN(n_5_1570));
   NAND2_X1 i_5_1306 (.A1(n_5_1569), .A2(n_5_1570), .ZN(n_5_1571));
   INV_X1 i_5_2030 (.A(m[11]), .ZN(n_5_1572));
   XNOR2_X1 i_5_2031 (.A(n_5_1749), .B(n_5_1367), .ZN(n_5_2007));
   NAND2_X1 i_5_2032 (.A1(n_5_3168), .A2(m[9]), .ZN(n_5_1573));
   INV_X1 i_5_2033 (.A(n_53), .ZN(n_5_1574));
   INV_X1 i_5_2034 (.A(n_54), .ZN(n_5_1575));
   INV_X1 i_5_2035 (.A(n_5_1816), .ZN(n_5_1576));
   INV_X1 i_5_2036 (.A(n_60), .ZN(n_5_1577));
   INV_X1 i_5_2037 (.A(n_73), .ZN(n_5_1578));
   INV_X1 i_5_2038 (.A(n_76), .ZN(n_5_1579));
   INV_X1 i_5_2039 (.A(n_75), .ZN(n_5_1580));
   INV_X1 i_5_2040 (.A(n_5_3191), .ZN(n_5_1581));
   INV_X1 i_5_2041 (.A(n_61), .ZN(n_5_1582));
   INV_X1 i_5_2042 (.A(n_5_3246), .ZN(n_5_1583));
   NAND2_X1 i_5_2043 (.A1(n_5_1583), .A2(n_5_1574), .ZN(n_5_1805));
   INV_X1 i_5_2044 (.A(n_5_1601), .ZN(n_5_1584));
   NAND2_X1 i_5_2045 (.A1(n_5_2924), .A2(n_5_1684), .ZN(n_5_1585));
   XNOR2_X1 i_5_2046 (.A(n_5_1812), .B(n_5_2568), .ZN(n_5_1586));
   XNOR2_X1 i_5_2047 (.A(n_5_1584), .B(n_5_1586), .ZN(n_5_1587));
   XNOR2_X1 i_5_2048 (.A(n_5_3107), .B(n_73), .ZN(n_5_1588));
   XNOR2_X1 i_5_2049 (.A(n_53), .B(n_5_1575), .ZN(n_5_1589));
   AND2_X1 i_5_2050 (.A1(n_5_1599), .A2(n_5_1623), .ZN(n_5_2214));
   INV_X1 i_5_2051 (.A(n_60), .ZN(n_5_1590));
   NAND2_X1 i_5_2052 (.A1(n_5_1611), .A2(n_5_1610), .ZN(n_5_1591));
   XOR2_X1 i_5_2053 (.A(n_5_2914), .B(n_5_1728), .Z(n_5_1592));
   OAI211_X1 i_5_1648 (.A(n_5_1706), .B(n_5_1614), .C1(n_5_1642), .C2(n_5_1668), 
      .ZN(n_5_1593));
   XOR2_X1 i_5_1322 (.A(n_5_1590), .B(n_5_1816), .Z(n_5_1594));
   NAND2_X1 i_5_2056 (.A1(n_5_1738), .A2(n_5_1741), .ZN(n_5_3178));
   NAND2_X1 i_5_2057 (.A1(n_5_1595), .A2(n_5_1636), .ZN(n_5_2216));
   NAND2_X1 i_5_2058 (.A1(n_5_1596), .A2(n_5_1671), .ZN(n_5_1595));
   NAND2_X1 i_5_2059 (.A1(n_5_1633), .A2(n_5_1613), .ZN(n_5_1596));
   INV_X1 i_5_2060 (.A(n_76), .ZN(n_5_1597));
   NAND2_X1 i_5_2061 (.A1(n_5_1667), .A2(n_5_1653), .ZN(n_5_1598));
   OAI21_X1 i_5_1323 (.A(n_5_1708), .B1(n_5_3733), .B2(n_5_2866), .ZN(n_5_1599));
   INV_X1 i_5_2063 (.A(n_5_3185), .ZN(n_5_1600));
   NAND2_X1 i_5_2064 (.A1(n_5_1811), .A2(m[0]), .ZN(n_5_1601));
   XNOR2_X1 i_5_2065 (.A(n_5_1661), .B(n_5_1651), .ZN(n_5_1602));
   NAND2_X1 i_5_2066 (.A1(n_5_1631), .A2(n_5_1605), .ZN(n_5_1603));
   NAND3_X1 i_5_2067 (.A1(n_5_1628), .A2(n_5_1677), .A3(n_5_1680), .ZN(n_5_1604));
   NAND4_X1 i_5_2068 (.A1(n_5_1644), .A2(n_5_1627), .A3(n_5_1700), .A4(n_5_1701), 
      .ZN(n_5_1605));
   INV_X1 i_5_2069 (.A(n_75), .ZN(n_5_1606));
   NAND2_X1 i_5_2070 (.A1(n_5_3187), .A2(n_5_1675), .ZN(n_5_2217));
   NOR2_X1 i_5_2071 (.A1(n_5_1812), .A2(n_5_2568), .ZN(n_5_1607));
   AOI22_X1 i_5_2072 (.A1(n_5_1812), .A2(n_5_2568), .B1(m[0]), .B2(n_5_1811), 
      .ZN(n_5_1608));
   INV_X1 i_5_2073 (.A(n_5_1610), .ZN(n_5_1609));
   NAND2_X1 i_5_2074 (.A1(n_5_3822), .A2(n_5_3329), .ZN(n_5_1610));
   OR2_X1 i_5_2075 (.A1(n_5_3822), .A2(n_5_3329), .ZN(n_5_1611));
   OAI21_X1 i_5_2076 (.A(n_5_1741), .B1(n_5_1740), .B2(n_5_1676), .ZN(n_5_1612));
   NAND2_X1 i_5_2077 (.A1(n_5_3111), .A2(n_5_1578), .ZN(n_5_1613));
   NAND2_X1 i_5_2078 (.A1(n_5_3554), .A2(n_66), .ZN(n_5_1614));
   NAND2_X1 i_5_2079 (.A1(n_5_1612), .A2(n_5_1613), .ZN(n_5_1615));
   NAND2_X1 i_5_2080 (.A1(n_5_2918), .A2(n_5_2569), .ZN(n_5_1616));
   NOR2_X1 i_5_2081 (.A1(n_5_2918), .A2(n_5_2569), .ZN(n_5_1617));
   NAND2_X1 i_5_2082 (.A1(n_5_3107), .A2(n_73), .ZN(n_5_1618));
   NAND2_X1 i_5_2083 (.A1(n_5_3107), .A2(n_73), .ZN(n_5_1619));
   INV_X1 i_5_2084 (.A(n_5_1619), .ZN(n_5_1620));
   XOR2_X1 i_5_2085 (.A(n_5_1670), .B(n_5_3548), .Z(n_5_1621));
   INV_X1 i_5_2086 (.A(n_5_1589), .ZN(n_5_2218));
   XNOR2_X1 i_5_2087 (.A(n_5_3342), .B(n_5_1675), .ZN(n_5_1622));
   OR2_X1 i_5_2088 (.A1(n_5_3733), .A2(n_5_2866), .ZN(n_5_2219));
   NAND2_X1 i_5_1325 (.A1(n_5_3733), .A2(n_5_2866), .ZN(n_5_1623));
   INV_X1 i_5_2090 (.A(n_5_2866), .ZN(n_5_1624));
   XNOR2_X1 i_5_1649 (.A(n_5_3733), .B(n_5_1624), .ZN(n_5_1625));
   INV_X1 i_5_1650 (.A(n_5_1593), .ZN(n_5_1626));
   NAND2_X1 i_5_2093 (.A1(n_5_1821), .A2(n_5_1606), .ZN(n_5_1627));
   NAND2_X1 i_5_2094 (.A1(n_5_4471), .A2(n_5_1579), .ZN(n_5_1628));
   NAND2_X1 i_5_2095 (.A1(n_5_4471), .A2(n_5_1579), .ZN(n_5_1629));
   INV_X1 i_5_2096 (.A(n_5_1615), .ZN(n_5_1630));
   NAND2_X1 i_5_2097 (.A1(n_5_1645), .A2(n_5_1604), .ZN(n_5_1631));
   NAND2_X1 i_5_2098 (.A1(n_5_1676), .A2(n_5_1741), .ZN(n_5_1632));
   NAND2_X1 i_5_2099 (.A1(n_5_1647), .A2(n_5_1618), .ZN(n_5_1633));
   INV_X1 i_5_2100 (.A(n_5_1613), .ZN(n_5_1634));
   AOI21_X1 i_5_2101 (.A(n_5_1634), .B1(n_5_1647), .B2(n_5_1618), .ZN(n_5_1635));
   NAND2_X1 i_5_2102 (.A1(n_5_1673), .A2(n_5_1635), .ZN(n_5_1636));
   INV_X1 i_5_1651 (.A(n_5_3412), .ZN(n_5_1637));
   INV_X1 i_5_2104 (.A(n_5_1624), .ZN(n_5_1638));
   XNOR2_X1 i_5_2105 (.A(n_5_1624), .B(n_5_1600), .ZN(n_5_1639));
   OAI22_X1 i_5_1653 (.A1(n_5_1637), .A2(n_5_1638), .B1(n_5_3412), .B2(n_5_1639), 
      .ZN(n_5_1640));
   INV_X1 i_5_2107 (.A(n_5_1738), .ZN(n_5_1641));
   NOR2_X1 i_5_2108 (.A1(n_5_3554), .A2(n_66), .ZN(n_5_1642));
   INV_X1 i_5_2109 (.A(n_5_1821), .ZN(n_5_1643));
   NAND2_X1 i_5_2110 (.A1(n_5_1643), .A2(n_75), .ZN(n_5_1644));
   AOI21_X1 i_5_2111 (.A(n_5_1690), .B1(n_5_1697), .B2(n_5_1648), .ZN(n_5_1645));
   INV_X1 i_5_2112 (.A(n_5_1741), .ZN(n_5_1646));
   OAI21_X1 i_5_2113 (.A(n_5_1632), .B1(n_5_1652), .B2(n_5_1646), .ZN(n_5_1647));
   NAND3_X1 i_5_2114 (.A1(n_5_1821), .A2(n_5_2962), .A3(n_5_1606), .ZN(n_5_1648));
   AOI21_X1 i_5_2115 (.A(n_5_1620), .B1(n_5_4462), .B2(n_76), .ZN(n_5_1649));
   NAND2_X1 i_5_2116 (.A1(n_5_1612), .A2(n_5_1613), .ZN(n_5_1650));
   AOI21_X1 i_5_2117 (.A(n_5_1642), .B1(n_5_1669), .B2(n_5_1614), .ZN(n_5_1651));
   NAND2_X1 i_5_2118 (.A1(n_5_1598), .A2(n_5_1740), .ZN(n_5_1652));
   NAND2_X1 i_5_2119 (.A1(n_5_1576), .A2(n_5_1577), .ZN(n_5_1653));
   INV_X1 i_5_2120 (.A(n_5_1740), .ZN(n_5_1654));
   NAND2_X1 i_5_2121 (.A1(n_5_1576), .A2(n_5_1577), .ZN(n_5_1655));
   NAND2_X1 i_5_2122 (.A1(n_5_1654), .A2(n_5_1655), .ZN(n_5_1656));
   INV_X1 i_5_2123 (.A(n_5_1655), .ZN(n_5_1657));
   OAI21_X1 i_5_2124 (.A(n_5_1656), .B1(n_5_1598), .B2(n_5_1657), .ZN(n_5_3179));
   INV_X1 i_5_2125 (.A(n_5_3412), .ZN(n_5_1658));
   INV_X1 i_5_2126 (.A(n_5_3185), .ZN(n_5_1659));
   INV_X1 i_5_2127 (.A(n_5_1600), .ZN(n_5_1660));
   OAI22_X1 i_5_2128 (.A1(n_5_1658), .A2(n_5_1659), .B1(n_5_3412), .B2(n_5_1660), 
      .ZN(n_5_1661));
   INV_X1 i_5_2129 (.A(n_61), .ZN(n_5_1662));
   XNOR2_X1 i_5_2130 (.A(n_5_3191), .B(n_5_1662), .ZN(n_5_1663));
   XNOR2_X1 i_5_2131 (.A(n_5_1756), .B(n_5_1663), .ZN(n_5_1664));
   NAND3_X1 i_5_1326 (.A1(n_5_1711), .A2(n_5_1599), .A3(n_5_1623), .ZN(n_5_1665));
   XNOR2_X1 i_5_1328 (.A(n_5_1594), .B(n_5_1665), .ZN(n_5_1666));
   NAND3_X1 i_5_2134 (.A1(n_5_1711), .A2(n_5_1599), .A3(n_5_1623), .ZN(n_5_1667));
   OAI21_X1 i_5_2135 (.A(n_5_3336), .B1(n_5_1674), .B2(n_5_3262), .ZN(n_5_1668));
   OAI21_X1 i_5_2136 (.A(n_5_3336), .B1(n_5_1674), .B2(n_5_3262), .ZN(n_5_1669));
   OAI21_X1 i_5_2137 (.A(n_5_3336), .B1(n_5_1674), .B2(n_5_3262), .ZN(n_5_1670));
   XNOR2_X1 i_5_2138 (.A(n_5_4462), .B(n_5_1597), .ZN(n_5_1671));
   INV_X1 i_5_2139 (.A(n_5_1597), .ZN(n_5_1672));
   XNOR2_X1 i_5_2140 (.A(n_5_4462), .B(n_5_1672), .ZN(n_5_1673));
   AOI21_X1 i_5_2141 (.A(n_5_1617), .B1(n_5_1729), .B2(n_5_1616), .ZN(n_5_1674));
   AOI21_X1 i_5_2142 (.A(n_5_1617), .B1(n_5_1728), .B2(n_5_1616), .ZN(n_5_1675));
   NOR2_X1 i_5_2143 (.A1(n_5_3094), .A2(n_55), .ZN(n_5_1676));
   NAND2_X1 i_5_2144 (.A1(n_5_2217), .A2(n_5_2214), .ZN(n_5_1677));
   INV_X1 i_5_2145 (.A(n_5_1641), .ZN(n_5_1678));
   NAND3_X1 i_5_2146 (.A1(n_5_1678), .A2(n_5_1613), .A3(n_5_1653), .ZN(n_5_1679));
   INV_X1 i_5_2147 (.A(n_5_1679), .ZN(n_5_1680));
   INV_X1 i_5_2148 (.A(n_53), .ZN(n_5_1681));
   XNOR2_X1 i_5_2149 (.A(n_5_3246), .B(n_5_1681), .ZN(n_5_1682));
   XNOR2_X1 i_5_2150 (.A(n_5_1585), .B(n_5_1682), .ZN(n_5_1683));
   NAND2_X1 i_5_2151 (.A1(n_5_1581), .A2(n_5_1582), .ZN(n_5_1684));
   NAND2_X1 i_5_2152 (.A1(n_5_1581), .A2(n_5_1582), .ZN(n_5_1685));
   NAND2_X1 i_5_2153 (.A1(n_5_1761), .A2(n_5_1685), .ZN(n_5_4066));
   NAND2_X1 i_5_2154 (.A1(n_5_1630), .A2(n_5_1629), .ZN(n_5_1686));
   NAND2_X1 i_5_2155 (.A1(n_5_3107), .A2(n_73), .ZN(n_5_1687));
   INV_X1 i_5_2156 (.A(n_5_1687), .ZN(n_5_1688));
   NAND2_X1 i_5_2157 (.A1(n_5_1628), .A2(n_5_1688), .ZN(n_5_1689));
   NAND2_X1 i_5_2158 (.A1(n_5_1686), .A2(n_5_1689), .ZN(n_5_1690));
   NAND2_X1 i_5_2159 (.A1(n_5_1675), .A2(n_5_3336), .ZN(n_5_1691));
   INV_X1 i_5_1330 (.A(n_5_1691), .ZN(n_5_1692));
   INV_X1 i_5_2161 (.A(n_5_2866), .ZN(n_5_1693));
   INV_X1 i_5_2162 (.A(n_5_1821), .ZN(n_5_1694));
   INV_X1 i_5_2163 (.A(n_75), .ZN(n_5_1695));
   AOI21_X1 i_5_2164 (.A(n_5_1695), .B1(n_5_4462), .B2(n_76), .ZN(n_5_1696));
   NAND2_X1 i_5_2165 (.A1(n_5_1694), .A2(n_5_1696), .ZN(n_5_1697));
   NAND2_X1 i_5_1847 (.A1(n_5_1626), .A2(n_5_1625), .ZN(n_5_1698));
   XNOR2_X1 i_5_1864 (.A(n_5_3733), .B(n_5_1640), .ZN(n_5_1699));
   OAI21_X1 i_5_1868 (.A(n_5_1698), .B1(n_5_1699), .B2(n_5_1626), .ZN(n_5_2221));
   NAND3_X1 i_5_2169 (.A1(n_5_1702), .A2(n_5_1649), .A3(n_5_1650), .ZN(n_5_1700));
   NAND3_X1 i_5_2170 (.A1(n_5_2962), .A2(n_5_4471), .A3(n_5_1579), .ZN(n_5_1701));
   NAND2_X1 i_5_2171 (.A1(n_5_1703), .A2(n_5_1704), .ZN(n_5_1702));
   INV_X1 i_5_2172 (.A(n_5_1752), .ZN(n_5_1703));
   NOR2_X1 i_5_2173 (.A1(n_5_1641), .A2(n_5_3104), .ZN(n_5_1704));
   NAND2_X1 i_5_2174 (.A1(n_5_1649), .A2(n_5_1650), .ZN(n_5_1705));
   NAND2_X1 i_5_2175 (.A1(n_5_3412), .A2(n_5_3185), .ZN(n_5_1706));
   NAND2_X1 i_5_2176 (.A1(n_5_3412), .A2(n_5_3185), .ZN(n_5_1707));
   NAND2_X1 i_5_1334 (.A1(n_5_1715), .A2(n_5_1707), .ZN(n_5_1708));
   INV_X1 i_5_2178 (.A(n_5_3733), .ZN(n_5_1709));
   NAND2_X1 i_5_1336 (.A1(n_5_1709), .A2(n_5_1693), .ZN(n_5_1710));
   NAND3_X1 i_5_1361 (.A1(n_5_3490), .A2(n_5_1710), .A3(n_5_1692), .ZN(n_5_1711));
   INV_X1 i_5_2181 (.A(n_5_3553), .ZN(n_5_3180));
   NAND2_X1 i_5_2182 (.A1(n_5_3414), .A2(n_5_1600), .ZN(n_5_3181));
   NAND2_X1 i_5_2183 (.A1(n_5_3554), .A2(n_66), .ZN(n_5_1712));
   AOI21_X1 i_5_2184 (.A(n_5_3549), .B1(n_5_3263), .B2(n_5_1712), .ZN(n_5_1713));
   INV_X1 i_5_2185 (.A(n_5_1600), .ZN(n_5_1714));
   OAI21_X1 i_5_2186 (.A(n_5_1713), .B1(n_5_3412), .B2(n_5_1714), .ZN(n_5_1715));
   NOR2_X1 i_5_2187 (.A1(n_5_2232), .A2(n_58), .ZN(n_5_1716));
   XNOR2_X1 i_5_2188 (.A(n_5_2232), .B(n_5_1285), .ZN(n_5_1717));
   XNOR2_X1 i_5_2189 (.A(n_5_2232), .B(m[4]), .ZN(n_5_1718));
   NAND3_X1 i_5_2190 (.A1(n_5_1456), .A2(n_5_1457), .A3(n_5_1436), .ZN(n_5_1719));
   NAND3_X1 i_5_2191 (.A1(n_5_2946), .A2(n_5_1454), .A3(n_5_1435), .ZN(n_5_1720));
   NAND2_X1 i_5_2192 (.A1(n_5_2012), .A2(n_5_2569), .ZN(n_5_1721));
   XNOR2_X1 i_5_2193 (.A(n_5_2012), .B(n_5_2569), .ZN(n_5_2225));
   NAND2_X1 i_5_2194 (.A1(n_5_2012), .A2(n_5_2569), .ZN(n_5_1722));
   INV_X1 i_5_2195 (.A(n_5_1720), .ZN(n_5_1723));
   INV_X1 i_5_2196 (.A(n_5_2012), .ZN(n_5_2010));
   NAND2_X1 i_5_2197 (.A1(n_5_1720), .A2(m[3]), .ZN(n_5_2011));
   XNOR2_X1 i_5_2198 (.A(n_5_1720), .B(n_5_1387), .ZN(n_5_1724));
   NAND3_X1 i_5_2199 (.A1(n_5_2946), .A2(n_5_1454), .A3(n_5_1435), .ZN(n_5_2012));
   XNOR2_X1 i_5_2200 (.A(n_5_1748), .B(n_5_1588), .ZN(n_5_1725));
   NAND2_X1 i_5_2201 (.A1(n_5_1725), .A2(n_5_1452), .ZN(n_5_1726));
   NOR2_X1 i_5_2202 (.A1(n_5_1608), .A2(n_5_1607), .ZN(n_5_1727));
   OAI21_X1 i_5_2203 (.A(n_5_1611), .B1(n_5_1727), .B2(n_5_1609), .ZN(n_5_1728));
   OAI21_X1 i_5_2204 (.A(n_5_1611), .B1(n_5_1730), .B2(n_5_1609), .ZN(n_5_1729));
   NOR2_X1 i_5_2205 (.A1(n_5_1608), .A2(n_5_1607), .ZN(n_5_1730));
   NAND2_X1 i_5_2206 (.A1(n_5_1446), .A2(n_5_1449), .ZN(n_5_1731));
   INV_X1 i_5_2207 (.A(n_5_1731), .ZN(n_5_1732));
   NAND2_X1 i_5_2208 (.A1(n_5_2013), .A2(m[12]), .ZN(n_5_1733));
   XNOR2_X1 i_5_2209 (.A(n_5_2013), .B(m[12]), .ZN(n_5_3182));
   XNOR2_X1 i_5_2210 (.A(n_5_1731), .B(n_75), .ZN(n_5_1734));
   NAND2_X1 i_5_2211 (.A1(n_5_1446), .A2(n_5_1449), .ZN(n_5_2013));
   NAND3_X1 i_5_2212 (.A1(n_5_2962), .A2(n_5_4471), .A3(n_5_1579), .ZN(n_5_1735));
   NAND3_X1 i_5_2213 (.A1(n_5_2962), .A2(n_5_4471), .A3(n_5_1579), .ZN(n_5_1736));
   NOR2_X1 i_5_2214 (.A1(n_5_1641), .A2(n_5_3104), .ZN(n_5_1737));
   INV_X1 i_5_2215 (.A(n_5_1739), .ZN(n_5_1738));
   NOR2_X1 i_5_2216 (.A1(n_5_3094), .A2(n_55), .ZN(n_5_1739));
   NAND2_X1 i_5_2217 (.A1(n_5_1816), .A2(n_60), .ZN(n_5_1740));
   NAND2_X1 i_5_2218 (.A1(n_5_3094), .A2(n_55), .ZN(n_5_1741));
   NAND2_X1 i_5_2219 (.A1(n_5_3094), .A2(n_55), .ZN(n_5_1742));
   NAND2_X1 i_5_2220 (.A1(n_5_1816), .A2(n_60), .ZN(n_5_1743));
   NAND2_X1 i_5_2221 (.A1(n_5_1742), .A2(n_5_1743), .ZN(n_5_1744));
   INV_X1 i_5_2222 (.A(n_5_1744), .ZN(n_5_1745));
   INV_X1 i_5_2223 (.A(n_5_1667), .ZN(n_5_1746));
   OAI21_X1 i_5_2224 (.A(n_5_1653), .B1(n_5_3094), .B2(n_55), .ZN(n_5_1747));
   AOI22_X1 i_5_2225 (.A1(n_5_1745), .A2(n_5_1746), .B1(n_5_1747), .B2(n_5_1742), 
      .ZN(n_5_1748));
   NAND2_X1 i_5_2226 (.A1(n_5_1455), .A2(n_5_1445), .ZN(n_5_2014));
   XNOR2_X1 i_5_2227 (.A(n_5_2014), .B(n_5_1572), .ZN(n_5_1749));
   OR2_X1 i_5_2228 (.A1(n_5_2014), .A2(n_76), .ZN(n_5_1750));
   NAND2_X1 i_5_2229 (.A1(n_5_1455), .A2(n_5_1445), .ZN(n_5_1751));
   NAND2_X1 i_5_2230 (.A1(n_5_1613), .A2(n_5_1653), .ZN(n_5_1752));
   NAND2_X1 i_5_2231 (.A1(n_5_1613), .A2(n_5_1653), .ZN(n_5_1753));
   INV_X1 i_5_2232 (.A(n_5_1753), .ZN(n_5_1754));
   NAND2_X1 i_5_2233 (.A1(n_5_3540), .A2(n_5_3133), .ZN(n_5_2228));
   INV_X1 i_5_2234 (.A(n_5_2228), .ZN(n_5_1755));
   AOI21_X1 i_5_2235 (.A(n_5_1808), .B1(n_5_3853), .B2(n_5_1810), .ZN(n_5_1756));
   INV_X1 i_5_2236 (.A(n_5_4195), .ZN(n_5_1808));
   NAND2_X1 i_5_2237 (.A1(n_5_1643), .A2(n_5_1580), .ZN(n_5_1810));
   NAND2_X1 i_5_2238 (.A1(n_5_1643), .A2(n_5_1580), .ZN(n_5_1757));
   INV_X1 i_5_2239 (.A(n_5_1757), .ZN(n_5_1758));
   NAND2_X1 i_5_2240 (.A1(n_5_4195), .A2(n_5_1758), .ZN(n_5_1759));
   NAND2_X1 i_5_2241 (.A1(n_5_4199), .A2(n_5_1759), .ZN(n_5_1760));
   INV_X1 i_5_2242 (.A(n_5_1760), .ZN(n_5_1761));
   NAND2_X1 i_5_2243 (.A1(n_5_3107), .A2(m[10]), .ZN(n_5_1762));
   NOR2_X1 i_5_2244 (.A1(n_5_3107), .A2(m[10]), .ZN(n_5_3183));
   XNOR2_X1 i_5_2245 (.A(n_5_3107), .B(m[10]), .ZN(n_5_1763));
   NAND2_X1 i_5_2246 (.A1(n_5_3243), .A2(n_5_3454), .ZN(n_5_1764));
   NAND2_X1 i_5_2247 (.A1(n_5_3222), .A2(n_5_1764), .ZN(n_5_1765));
   NAND2_X1 i_5_2248 (.A1(n_5_1683), .A2(n_5_1452), .ZN(n_5_1766));
   NAND2_X1 i_5_2249 (.A1(n_5_3216), .A2(n_5_3170), .ZN(n_5_1767));
   NAND2_X1 i_5_2250 (.A1(n_5_3216), .A2(n_5_3170), .ZN(n_5_1768));
   INV_X1 i_5_2251 (.A(n_5_3171), .ZN(n_5_1769));
   AOI21_X1 i_5_2252 (.A(n_5_1769), .B1(n_5_1683), .B2(n_5_1452), .ZN(n_5_1770));
   NAND2_X1 i_5_2253 (.A1(n_5_1768), .A2(n_5_1770), .ZN(n_5_2017));
   INV_X1 i_5_2254 (.A(n_5_3162), .ZN(n_5_2229));
   NAND2_X1 i_5_2255 (.A1(n_5_1479), .A2(n_5_1525), .ZN(n_5_1771));
   NAND2_X1 i_5_2256 (.A1(n_5_1479), .A2(n_5_1525), .ZN(n_5_1772));
   AOI21_X1 i_5_2257 (.A(n_5_3550), .B1(n_5_1772), .B2(n_5_3551), .ZN(n_5_1773));
   AOI21_X1 i_5_2258 (.A(n_5_3550), .B1(n_5_1771), .B2(n_5_3551), .ZN(n_5_1774));
   XOR2_X1 i_5_2259 (.A(n_5_1772), .B(n_5_3552), .Z(n_5_1775));
   NAND3_X1 i_5_2260 (.A1(n_5_1273), .A2(n_5_1281), .A3(n_5_1750), .ZN(n_5_1776));
   NAND2_X1 i_5_2261 (.A1(n_5_1751), .A2(n_76), .ZN(n_5_1777));
   NAND2_X1 i_5_2262 (.A1(n_5_1776), .A2(n_5_1777), .ZN(n_5_1778));
   NAND2_X1 i_5_2263 (.A1(n_5_1561), .A2(m[13]), .ZN(n_5_1779));
   INV_X1 i_5_2264 (.A(n_5_1347), .ZN(n_5_1780));
   NAND2_X1 i_5_2265 (.A1(n_5_1561), .A2(m[13]), .ZN(n_5_1781));
   NAND2_X1 i_5_2266 (.A1(n_5_1780), .A2(n_5_1781), .ZN(n_5_1782));
   XNOR2_X1 i_5_2267 (.A(n_5_3261), .B(m[6]), .ZN(n_5_1783));
   NAND3_X1 i_5_2268 (.A1(n_5_1437), .A2(n_5_1438), .A3(n_5_1439), .ZN(n_5_1784));
   NAND2_X1 i_5_2269 (.A1(n_5_1300), .A2(n_5_1327), .ZN(n_5_1785));
   NAND2_X1 i_5_2270 (.A1(n_5_1723), .A2(n_5_1301), .ZN(n_5_1786));
   NAND2_X1 i_5_2271 (.A1(n_5_1300), .A2(n_5_1327), .ZN(n_5_1787));
   NAND2_X1 i_5_2272 (.A1(n_5_1723), .A2(n_5_1301), .ZN(n_5_1790));
   XNOR2_X1 i_5_2273 (.A(n_5_3102), .B(n_5_1763), .ZN(n_5_1788));
   NAND2_X1 i_5_2274 (.A1(n_5_1788), .A2(n_5_3170), .ZN(n_5_1789));
   NAND2_X1 i_5_2275 (.A1(n_5_1719), .A2(n_58), .ZN(n_5_1791));
   NAND2_X1 i_5_2276 (.A1(n_5_1719), .A2(n_58), .ZN(n_5_1792));
   INV_X1 i_5_2277 (.A(n_5_1792), .ZN(n_5_2022));
   NAND3_X1 i_5_2278 (.A1(n_5_1456), .A2(n_5_1457), .A3(n_5_1436), .ZN(n_5_2232));
   NAND3_X1 i_5_2279 (.A1(n_5_1457), .A2(n_5_1456), .A3(n_5_1436), .ZN(n_5_2233));
   NAND3_X1 i_5_2280 (.A1(n_5_1437), .A2(n_5_1438), .A3(n_5_1439), .ZN(n_5_2234));
   OAI21_X1 i_5_2281 (.A(n_5_2187), .B1(n_5_2188), .B2(n_5_2211), .ZN(n_5_2025));
   NAND2_X1 i_5_2282 (.A1(n_5_3096), .A2(n_5_1461), .ZN(n_5_2235));
   INV_X1 i_5_2283 (.A(n_5_1481), .ZN(n_5_2236));
   NAND2_X1 i_5_2284 (.A1(n_5_3096), .A2(n_5_1461), .ZN(n_5_2237));
   NAND2_X1 i_5_2285 (.A1(n_5_1857), .A2(n_5_4069), .ZN(n_5_1793));
   NAND2_X1 i_5_2286 (.A1(n_5_2120), .A2(n_5_4068), .ZN(n_5_1794));
   NAND2_X1 i_5_2287 (.A1(n_5_1824), .A2(n_5_2886), .ZN(n_5_1795));
   NAND3_X1 i_5_2288 (.A1(n_5_1793), .A2(n_5_1794), .A3(n_5_1795), .ZN(n_5_1811));
   NAND2_X1 i_5_2289 (.A1(n_5_1859), .A2(n_5_4069), .ZN(n_5_1796));
   NAND2_X1 i_5_2290 (.A1(n_5_2177), .A2(n_5_4068), .ZN(n_5_1797));
   NAND2_X1 i_5_2291 (.A1(n_5_1824), .A2(n_5_2867), .ZN(n_5_1798));
   NAND3_X1 i_5_2292 (.A1(n_5_1796), .A2(n_5_1797), .A3(n_5_1798), .ZN(n_5_1812));
   NAND2_X1 i_5_2293 (.A1(n_5_2795), .A2(n_5_1824), .ZN(n_5_1799));
   NAND2_X1 i_5_2294 (.A1(n_5_2812), .A2(n_5_1824), .ZN(n_5_1813));
   NAND2_X1 i_5_2295 (.A1(n_5_2803), .A2(n_5_1824), .ZN(n_5_2238));
   NAND2_X1 i_5_2296 (.A1(n_5_2824), .A2(n_5_1824), .ZN(n_5_1800));
   NAND2_X1 i_5_2297 (.A1(n_5_2570), .A2(n_5_1824), .ZN(n_5_2239));
   NAND2_X1 i_5_2298 (.A1(n_5_2896), .A2(n_5_1824), .ZN(n_5_1801));
   INV_X1 i_5_2299 (.A(n_5_1801), .ZN(n_5_3389));
   NAND2_X1 i_5_1463 (.A1(n_5_3130), .A2(n_5_1824), .ZN(n_5_1802));
   INV_X1 i_5_1482 (.A(n_5_1802), .ZN(n_5_1807));
   AOI21_X1 i_5_1483 (.A(n_5_1807), .B1(n_5_2070), .B2(n_5_4069), .ZN(n_5_1809));
   NAND2_X1 i_5_1515 (.A1(n_5_3078), .A2(n_5_1809), .ZN(n_5_1816));
   NAND2_X1 i_5_2304 (.A1(n_5_2336), .A2(n_5_1824), .ZN(n_5_2240));
   NAND2_X1 i_5_2305 (.A1(n_5_2292), .A2(n_5_4068), .ZN(n_5_2241));
   NAND2_X1 i_5_2306 (.A1(n_5_1870), .A2(n_5_4069), .ZN(n_5_2242));
   NAND2_X1 i_5_2307 (.A1(n_5_2340), .A2(n_5_1824), .ZN(n_5_2243));
   NAND2_X1 i_5_2308 (.A1(n_5_2344), .A2(n_5_1824), .ZN(n_5_4067));
   NAND2_X1 i_5_2309 (.A1(n_5_2115), .A2(n_5_4068), .ZN(n_5_1814));
   NAND2_X1 i_5_2310 (.A1(n_5_1879), .A2(n_5_4069), .ZN(n_5_1815));
   NAND2_X1 i_5_2311 (.A1(n_5_2347), .A2(n_5_1824), .ZN(n_5_1818));
   NAND3_X1 i_5_2312 (.A1(n_5_1814), .A2(n_5_1815), .A3(n_5_1818), .ZN(n_5_1821));
   INV_X1 i_5_2313 (.A(r[1]), .ZN(n_5_1822));
   NAND2_X1 i_5_2314 (.A1(r[2]), .A2(n_5_1822), .ZN(n_5_1823));
   INV_X1 i_5_2315 (.A(n_5_1823), .ZN(n_5_4068));
   NAND2_X1 i_5_2316 (.A1(n_5_2119), .A2(n_5_4068), .ZN(n_5_2245));
   NOR2_X1 i_5_2317 (.A1(r[2]), .A2(n_5_1822), .ZN(n_5_4069));
   NAND2_X1 i_5_2318 (.A1(n_5_1856), .A2(n_5_4069), .ZN(n_5_2247));
   XNOR2_X1 i_5_2319 (.A(r[2]), .B(r[1]), .ZN(n_5_1824));
   NAND2_X1 i_5_2320 (.A1(n_5_2354), .A2(n_5_1824), .ZN(n_5_2248));
   NAND2_X1 i_5_2321 (.A1(n_5_2175), .A2(n_5_4068), .ZN(n_5_1825));
   NAND2_X1 i_5_2322 (.A1(n_5_1865), .A2(n_5_4069), .ZN(n_5_1827));
   NAND2_X1 i_5_2323 (.A1(n_5_2222), .A2(n_5_4068), .ZN(n_5_1829));
   NAND2_X1 i_5_2324 (.A1(n_5_1862), .A2(n_5_4069), .ZN(n_5_1830));
   NAND2_X1 i_5_2325 (.A1(n_5_2123), .A2(n_5_4068), .ZN(n_5_2249));
   NAND2_X1 i_5_2326 (.A1(n_5_2026), .A2(n_5_4069), .ZN(n_5_2250));
   NAND2_X1 i_5_2327 (.A1(n_5_2128), .A2(n_5_4068), .ZN(n_5_2251));
   NAND2_X1 i_5_2328 (.A1(n_5_1868), .A2(n_5_4069), .ZN(n_5_2252));
   NAND2_X1 i_5_2329 (.A1(n_5_2047), .A2(n_5_4069), .ZN(n_5_1831));
   NAND2_X1 i_5_2330 (.A1(n_5_2273), .A2(n_5_4068), .ZN(n_5_1832));
   INV_X1 i_5_2331 (.A(m[14]), .ZN(n_5_1833));
   INV_X1 i_5_2332 (.A(m[15]), .ZN(n_5_1834));
   INV_X1 i_5_2333 (.A(n_5_2344), .ZN(n_5_1835));
   INV_X1 i_5_2334 (.A(m[12]), .ZN(n_5_1836));
   INV_X1 i_5_2335 (.A(n_5_2347), .ZN(n_5_1837));
   INV_X1 i_5_2336 (.A(m[13]), .ZN(n_5_1838));
   NAND2_X1 i_5_2337 (.A1(n_5_1837), .A2(n_5_1838), .ZN(n_5_1839));
   NAND2_X1 i_5_2338 (.A1(n_5_2347), .A2(m[13]), .ZN(n_5_1840));
   NAND2_X1 i_5_2339 (.A1(n_5_2354), .A2(m[14]), .ZN(n_5_1841));
   INV_X1 i_5_2340 (.A(n_5_2354), .ZN(n_5_1842));
   NAND2_X1 i_5_2341 (.A1(n_5_1842), .A2(n_5_1833), .ZN(n_5_1843));
   INV_X1 i_5_2342 (.A(n_5_1840), .ZN(n_5_1845));
   INV_X1 i_5_2343 (.A(n_5_1891), .ZN(n_5_1846));
   INV_X1 i_5_2344 (.A(n_5_2055), .ZN(n_5_1847));
   AOI21_X1 i_5_2345 (.A(n_5_1846), .B1(n_5_1847), .B2(n_5_1885), .ZN(n_5_1848));
   NAND2_X1 i_5_2346 (.A1(n_5_2055), .A2(n_5_1891), .ZN(n_5_1849));
   NAND3_X1 i_5_2347 (.A1(n_5_1840), .A2(n_5_1849), .A3(n_5_1885), .ZN(n_5_1851));
   NAND3_X1 i_5_2348 (.A1(n_5_1851), .A2(n_5_1841), .A3(n_5_1839), .ZN(n_5_1852));
   NAND2_X1 i_5_2349 (.A1(n_5_1852), .A2(n_5_1843), .ZN(n_5_1853));
   XNOR2_X1 i_5_2350 (.A(n_5_2354), .B(m[14]), .ZN(n_5_1854));
   XNOR2_X1 i_5_2351 (.A(n_5_2815), .B(n_5_1854), .ZN(n_5_2253));
   XNOR2_X1 i_5_2352 (.A(m[14]), .B(n_5_1834), .ZN(n_5_1855));
   XNOR2_X1 i_5_2353 (.A(n_5_1853), .B(n_5_1855), .ZN(n_5_1856));
   XOR2_X1 i_5_2354 (.A(n_5_1940), .B(n_5_1858), .Z(n_5_1857));
   NAND2_X1 i_5_2355 (.A1(n_5_2865), .A2(m[0]), .ZN(n_5_1858));
   XNOR2_X1 i_5_2356 (.A(n_5_1861), .B(n_5_1860), .ZN(n_5_1859));
   NAND2_X1 i_5_2357 (.A1(n_5_2075), .A2(n_5_2805), .ZN(n_5_1860));
   NOR2_X1 i_5_2358 (.A1(n_5_2830), .A2(n_5_1935), .ZN(n_5_1861));
   XNOR2_X1 i_5_2359 (.A(n_5_1864), .B(n_5_1909), .ZN(n_5_1862));
   NOR2_X1 i_5_2360 (.A1(n_5_1896), .A2(n_5_2040), .ZN(n_5_1864));
   XNOR2_X1 i_5_2361 (.A(n_5_1910), .B(n_5_1866), .ZN(n_5_1865));
   NAND2_X1 i_5_2362 (.A1(n_5_1933), .A2(n_5_1921), .ZN(n_5_1866));
   XNOR2_X1 i_5_2363 (.A(n_5_2261), .B(n_5_1867), .ZN(n_5_3392));
   NAND2_X1 i_5_2364 (.A1(n_5_2027), .A2(n_5_2030), .ZN(n_5_1867));
   XNOR2_X1 i_5_2365 (.A(n_5_1900), .B(n_5_1869), .ZN(n_5_1868));
   AOI21_X1 i_5_2366 (.A(n_5_1906), .B1(n_5_2065), .B2(n_5_2033), .ZN(n_5_1869));
   NAND2_X1 i_5_2367 (.A1(n_5_1872), .A2(n_5_1875), .ZN(n_5_1870));
   NAND2_X1 i_5_2368 (.A1(n_5_1873), .A2(n_5_1874), .ZN(n_5_1872));
   NOR2_X1 i_5_2369 (.A1(n_5_1876), .A2(n_5_1899), .ZN(n_5_1873));
   NAND2_X1 i_5_2370 (.A1(n_5_2255), .A2(n_5_1887), .ZN(n_5_1874));
   OAI211_X1 i_5_2371 (.A(n_5_2255), .B(n_5_1887), .C1(n_5_1876), .C2(n_5_1899), 
      .ZN(n_5_1875));
   AOI21_X1 i_5_2372 (.A(n_5_1877), .B1(n_5_1878), .B2(n_5_2254), .ZN(n_5_1876));
   NAND2_X1 i_5_2373 (.A1(n_5_1898), .A2(n_5_2033), .ZN(n_5_1877));
   NAND3_X1 i_5_2374 (.A1(n_5_2071), .A2(n_5_2027), .A3(n_5_2072), .ZN(n_5_1878));
   NAND2_X1 i_5_2375 (.A1(n_5_1880), .A2(n_5_1882), .ZN(n_5_1879));
   NAND2_X1 i_5_2376 (.A1(n_5_1881), .A2(n_5_1901), .ZN(n_5_1880));
   NAND2_X1 i_5_2377 (.A1(n_5_1884), .A2(n_5_1891), .ZN(n_5_1881));
   NAND3_X1 i_5_2378 (.A1(n_5_1884), .A2(n_5_1891), .A3(n_5_1903), .ZN(n_5_1882));
   INV_X1 i_5_2379 (.A(m[13]), .ZN(n_5_1883));
   NAND3_X1 i_5_2380 (.A1(n_5_2041), .A2(n_5_2042), .A3(n_5_1885), .ZN(n_5_1884));
   NAND2_X1 i_5_2381 (.A1(n_5_2344), .A2(m[12]), .ZN(n_5_1885));
   NAND3_X1 i_5_2382 (.A1(n_5_1888), .A2(n_5_1887), .A3(n_5_1898), .ZN(n_5_1886));
   NAND2_X1 i_5_2383 (.A1(n_5_2340), .A2(m[11]), .ZN(n_5_1887));
   NAND2_X1 i_5_2384 (.A1(n_5_2256), .A2(n_5_1889), .ZN(n_5_1888));
   AOI21_X1 i_5_2385 (.A(n_5_1906), .B1(n_5_2027), .B2(n_5_2033), .ZN(n_5_1889));
   AOI21_X1 i_5_2386 (.A(n_5_1906), .B1(n_5_1890), .B2(n_5_2900), .ZN(n_5_2254));
   INV_X1 i_5_2387 (.A(m[8]), .ZN(n_5_1890));
   OR2_X1 i_5_2388 (.A1(n_5_2340), .A2(m[11]), .ZN(n_5_2255));
   NAND2_X1 i_5_2389 (.A1(n_5_1835), .A2(n_5_1836), .ZN(n_5_1891));
   INV_X1 i_5_2390 (.A(m[3]), .ZN(n_5_1892));
   INV_X1 i_5_2391 (.A(m[0]), .ZN(n_5_1893));
   OAI21_X1 i_5_2392 (.A(n_5_1894), .B1(n_5_1905), .B2(n_5_1895), .ZN(n_5_4070));
   NAND3_X1 i_5_2393 (.A1(n_5_1895), .A2(n_5_2042), .A3(n_5_2041), .ZN(n_5_1894));
   XOR2_X1 i_5_2394 (.A(m[12]), .B(n_5_2344), .Z(n_5_1895));
   AOI21_X1 i_5_2395 (.A(n_5_2037), .B1(n_5_1908), .B2(n_5_2075), .ZN(n_5_1896));
   INV_X1 i_5_2396 (.A(m[3]), .ZN(n_5_1897));
   INV_X1 i_5_2397 (.A(n_5_1899), .ZN(n_5_2256));
   NAND2_X1 i_5_2398 (.A1(n_5_2336), .A2(m[10]), .ZN(n_5_1898));
   NOR2_X1 i_5_2399 (.A1(n_5_2336), .A2(m[10]), .ZN(n_5_1899));
   XNOR2_X1 i_5_2400 (.A(n_5_2336), .B(m[10]), .ZN(n_5_1900));
   XNOR2_X1 i_5_2401 (.A(n_5_2347), .B(n_5_1883), .ZN(n_5_1901));
   INV_X1 i_5_2402 (.A(n_5_1883), .ZN(n_5_1902));
   XNOR2_X1 i_5_2403 (.A(n_5_2347), .B(n_5_1902), .ZN(n_5_1903));
   NAND2_X1 i_5_2404 (.A1(n_5_2042), .A2(n_5_2041), .ZN(n_5_1904));
   INV_X1 i_5_2405 (.A(n_5_1904), .ZN(n_5_1905));
   NOR2_X1 i_5_2406 (.A1(n_5_3130), .A2(m[9]), .ZN(n_5_1906));
   INV_X1 i_5_2407 (.A(m[9]), .ZN(n_5_1907));
   OAI21_X1 i_5_2408 (.A(n_5_2805), .B1(n_5_2830), .B2(n_5_1935), .ZN(n_5_1908));
   XNOR2_X1 i_5_2409 (.A(n_5_2812), .B(m[4]), .ZN(n_5_1909));
   NOR2_X1 i_5_2410 (.A1(n_5_1955), .A2(n_5_2797), .ZN(n_5_1910));
   NOR2_X1 i_5_2411 (.A1(n_5_2790), .A2(n_5_2009), .ZN(n_5_1911));
   INV_X1 i_5_2412 (.A(n_5_2812), .ZN(n_5_1912));
   INV_X1 i_5_2413 (.A(m[4]), .ZN(n_5_1913));
   NAND2_X1 i_5_2414 (.A1(n_5_2865), .A2(m[0]), .ZN(n_5_1914));
   NAND3_X1 i_5_2415 (.A1(n_5_2886), .A2(n_5_2865), .A3(m[0]), .ZN(n_5_1915));
   NAND2_X1 i_5_2416 (.A1(n_5_2867), .A2(m[2]), .ZN(n_5_1916));
   NAND2_X1 i_5_2417 (.A1(m[0]), .A2(m[1]), .ZN(n_5_1917));
   INV_X1 i_5_2418 (.A(n_5_1917), .ZN(n_5_1918));
   NAND2_X1 i_5_2419 (.A1(n_5_2865), .A2(n_5_1918), .ZN(n_5_1919));
   NAND2_X1 i_5_2420 (.A1(n_5_2795), .A2(m[3]), .ZN(n_5_1920));
   NAND2_X1 i_5_2421 (.A1(n_5_2824), .A2(m[6]), .ZN(n_5_1921));
   INV_X1 i_5_2422 (.A(m[6]), .ZN(n_5_1922));
   INV_X1 i_5_2423 (.A(m[5]), .ZN(n_5_1925));
   NAND2_X1 i_5_2424 (.A1(n_5_1922), .A2(n_5_1925), .ZN(n_5_1926));
   NAND2_X1 i_5_2425 (.A1(n_5_2886), .A2(m[1]), .ZN(n_5_1927));
   NAND2_X1 i_5_2426 (.A1(n_5_2886), .A2(m[1]), .ZN(n_5_1928));
   NAND2_X1 i_5_2427 (.A1(n_5_2889), .A2(n_5_1921), .ZN(n_5_1929));
   INV_X1 i_5_2428 (.A(n_5_2824), .ZN(n_5_1930));
   INV_X1 i_5_2429 (.A(m[6]), .ZN(n_5_1931));
   NAND2_X1 i_5_2430 (.A1(n_5_1930), .A2(n_5_1931), .ZN(n_5_1932));
   OR2_X1 i_5_2431 (.A1(n_5_2824), .A2(m[6]), .ZN(n_5_1933));
   NAND2_X1 i_5_2432 (.A1(n_5_2803), .A2(m[5]), .ZN(n_5_1934));
   NOR2_X1 i_5_2433 (.A1(n_5_2886), .A2(m[1]), .ZN(n_5_1935));
   INV_X1 i_5_2434 (.A(n_5_2886), .ZN(n_5_1936));
   INV_X1 i_5_2435 (.A(m[1]), .ZN(n_5_1937));
   NAND2_X1 i_5_2436 (.A1(n_5_1936), .A2(n_5_1937), .ZN(n_5_1939));
   NAND2_X1 i_5_2437 (.A1(n_5_1939), .A2(n_5_1928), .ZN(n_5_1940));
   NAND2_X1 i_5_2438 (.A1(n_5_2812), .A2(m[4]), .ZN(n_5_1941));
   NAND3_X1 i_5_2439 (.A1(n_5_2039), .A2(n_5_2810), .A3(n_5_2799), .ZN(n_5_1948));
   NAND3_X1 i_5_2440 (.A1(n_5_2080), .A2(n_5_2039), .A3(n_5_1941), .ZN(n_5_1949));
   AOI21_X1 i_5_2441 (.A(n_5_1961), .B1(n_5_1949), .B2(n_5_2015), .ZN(n_5_1955));
   NAND3_X1 i_5_2442 (.A1(n_5_2080), .A2(n_5_2039), .A3(n_5_1941), .ZN(n_5_1957));
   INV_X1 i_5_2443 (.A(n_5_1963), .ZN(n_5_1961));
   NAND2_X1 i_5_2444 (.A1(n_5_2803), .A2(m[5]), .ZN(n_5_1963));
   INV_X1 i_5_2445 (.A(m[5]), .ZN(n_5_1965));
   NAND2_X1 i_5_2446 (.A1(n_5_2037), .A2(n_5_2076), .ZN(n_5_2257));
   NAND2_X1 i_5_2447 (.A1(n_5_1926), .A2(m[6]), .ZN(n_5_2258));
   OAI21_X1 i_5_2448 (.A(n_5_3252), .B1(n_5_2824), .B2(n_5_1948), .ZN(n_5_1975));
   OAI21_X1 i_5_2449 (.A(n_5_3252), .B1(n_5_1948), .B2(n_5_2824), .ZN(n_5_1985));
   NAND3_X1 i_5_2450 (.A1(n_5_2076), .A2(n_5_2075), .A3(n_5_2074), .ZN(n_5_1990));
   NAND2_X1 i_5_2451 (.A1(n_5_1985), .A2(n_5_1990), .ZN(n_5_1991));
   NAND2_X1 i_5_2452 (.A1(n_5_1914), .A2(n_5_1927), .ZN(n_5_1992));
   INV_X1 i_5_2453 (.A(n_5_1992), .ZN(n_5_1993));
   OAI21_X1 i_5_2454 (.A(n_5_2805), .B1(n_5_1993), .B2(n_5_1935), .ZN(n_5_1994));
   NAND3_X1 i_5_2455 (.A1(n_5_1991), .A2(n_5_1929), .A3(n_5_1932), .ZN(n_5_2259));
   NAND2_X1 i_5_2456 (.A1(n_5_3226), .A2(n_5_2072), .ZN(n_5_1995));
   INV_X1 i_5_2457 (.A(n_5_1995), .ZN(n_5_2260));
   NOR2_X1 i_5_2458 (.A1(n_5_2867), .A2(m[2]), .ZN(n_5_2009));
   OR2_X1 i_5_2459 (.A1(n_5_2812), .A2(m[4]), .ZN(n_5_2015));
   INV_X1 i_5_2460 (.A(n_5_1957), .ZN(n_5_2018));
   NAND2_X1 i_5_2461 (.A1(n_5_2018), .A2(n_5_2798), .ZN(n_5_2019));
   XNOR2_X1 i_5_2462 (.A(n_5_1965), .B(m[4]), .ZN(n_5_2020));
   MUX2_X1 i_5_2463 (.A(n_5_2801), .B(n_5_2798), .S(n_5_2812), .Z(n_5_2021));
   OAI21_X1 i_5_2464 (.A(n_5_2019), .B1(n_5_2021), .B2(n_5_2018), .ZN(n_5_2026));
   NAND2_X1 i_5_2465 (.A1(n_5_2896), .A2(m[8]), .ZN(n_5_2027));
   NAND2_X1 i_5_2466 (.A1(n_5_2900), .A2(n_5_1890), .ZN(n_5_2030));
   NAND2_X1 i_5_2467 (.A1(n_5_3130), .A2(m[9]), .ZN(n_5_2033));
   INV_X1 i_5_2468 (.A(m[9]), .ZN(n_5_2034));
   INV_X1 i_5_2469 (.A(n_5_1907), .ZN(n_5_2035));
   NAND2_X1 i_5_2470 (.A1(n_5_1845), .A2(n_5_1839), .ZN(n_5_2036));
   INV_X1 i_5_2471 (.A(n_5_2789), .ZN(n_5_2037));
   INV_X1 i_5_2472 (.A(n_5_2795), .ZN(n_5_2038));
   NAND2_X1 i_5_2473 (.A1(n_5_2795), .A2(m[3]), .ZN(n_5_2039));
   NOR2_X1 i_5_2474 (.A1(n_5_2795), .A2(m[3]), .ZN(n_5_2040));
   NAND2_X1 i_5_2475 (.A1(n_5_3156), .A2(n_5_2261), .ZN(n_5_2041));
   NAND2_X1 i_5_2476 (.A1(n_5_1886), .A2(n_5_2255), .ZN(n_5_2042));
   NAND2_X1 i_5_2477 (.A1(n_5_2896), .A2(m[8]), .ZN(n_5_2043));
   NAND3_X1 i_5_2478 (.A1(n_5_2062), .A2(n_5_2063), .A3(n_5_2061), .ZN(n_5_2044));
   NAND2_X1 i_5_2479 (.A1(n_5_2570), .A2(m[7]), .ZN(n_5_2045));
   NAND2_X1 i_5_2480 (.A1(n_5_1911), .A2(n_5_1994), .ZN(n_5_2046));
   OAI21_X1 i_5_2481 (.A(n_5_2046), .B1(n_5_2048), .B2(n_5_2791), .ZN(n_5_2047));
   OAI21_X1 i_5_2482 (.A(n_5_1920), .B1(n_5_2060), .B2(n_5_2009), .ZN(n_5_2048));
   NAND3_X1 i_5_1516 (.A1(n_5_2044), .A2(n_5_2043), .A3(n_5_2045), .ZN(n_5_2052));
   NAND2_X1 i_5_1570 (.A1(n_5_2900), .A2(n_5_1890), .ZN(n_5_2053));
   NAND2_X1 i_5_2485 (.A1(n_5_1886), .A2(n_5_2255), .ZN(n_5_2054));
   NAND2_X1 i_5_2486 (.A1(n_5_3169), .A2(n_5_2054), .ZN(n_5_2055));
   INV_X1 i_5_2487 (.A(n_5_1893), .ZN(n_5_2056));
   NAND2_X1 i_5_2488 (.A1(n_5_2865), .A2(n_5_2056), .ZN(n_5_2057));
   NOR2_X1 i_5_2489 (.A1(n_5_1935), .A2(n_5_2057), .ZN(n_5_2058));
   NAND2_X1 i_5_2490 (.A1(n_5_2805), .A2(n_5_1928), .ZN(n_5_2059));
   NOR2_X1 i_5_2491 (.A1(n_5_2058), .A2(n_5_2059), .ZN(n_5_2060));
   NOR2_X1 i_5_2492 (.A1(n_5_3223), .A2(n_5_2831), .ZN(n_5_2061));
   NAND2_X1 i_5_2493 (.A1(n_5_1975), .A2(n_5_2080), .ZN(n_5_2062));
   NAND2_X1 i_5_2494 (.A1(n_5_2889), .A2(n_5_1921), .ZN(n_5_2063));
   INV_X1 i_5_2495 (.A(m[2]), .ZN(n_5_2064));
   NAND2_X1 i_5_2496 (.A1(n_5_2052), .A2(n_5_2053), .ZN(n_5_2065));
   INV_X1 i_5_1571 (.A(n_5_2052), .ZN(n_5_2066));
   NAND2_X1 i_5_2498 (.A1(n_5_2034), .A2(n_5_2035), .ZN(n_5_2067));
   NAND2_X1 i_5_1608 (.A1(n_5_2066), .A2(n_5_3033), .ZN(n_5_2068));
   XNOR2_X1 i_5_1609 (.A(n_5_3033), .B(n_5_2053), .ZN(n_5_2069));
   OAI21_X1 i_5_1610 (.A(n_5_2068), .B1(n_5_2069), .B2(n_5_2066), .ZN(n_5_2070));
   NAND3_X1 i_5_2502 (.A1(n_5_2879), .A2(n_5_2878), .A3(n_5_2877), .ZN(n_5_2071));
   NAND2_X1 i_5_2503 (.A1(n_5_2570), .A2(m[7]), .ZN(n_5_2072));
   NAND2_X1 i_5_2504 (.A1(n_5_2570), .A2(m[7]), .ZN(n_5_2073));
   NAND2_X1 i_5_2505 (.A1(n_5_2883), .A2(n_5_2073), .ZN(n_5_2261));
   NAND4_X1 i_5_2506 (.A1(n_5_1915), .A2(n_5_1916), .A3(n_5_1928), .A4(n_5_1919), 
      .ZN(n_5_2074));
   NAND2_X1 i_5_2507 (.A1(n_5_2873), .A2(n_5_2064), .ZN(n_5_2075));
   NAND2_X1 i_5_2508 (.A1(n_5_2038), .A2(n_5_1897), .ZN(n_5_2076));
   NAND4_X1 i_5_2509 (.A1(n_5_1916), .A2(n_5_1928), .A3(n_5_1915), .A4(n_5_1919), 
      .ZN(n_5_2077));
   NAND2_X1 i_5_2510 (.A1(n_5_2038), .A2(n_5_1897), .ZN(n_5_2078));
   NAND2_X1 i_5_2511 (.A1(n_5_2873), .A2(n_5_2064), .ZN(n_5_2079));
   NAND3_X1 i_5_2512 (.A1(n_5_2077), .A2(n_5_2078), .A3(n_5_2079), .ZN(n_5_2080));
   INV_X1 i_5_2513 (.A(n_53), .ZN(n_5_2081));
   INV_X1 i_5_2514 (.A(n_54), .ZN(n_5_2082));
   INV_X1 i_5_2515 (.A(n_5_2896), .ZN(n_5_2083));
   INV_X1 i_5_2516 (.A(n_60), .ZN(n_5_2084));
   INV_X1 i_5_2517 (.A(n_5_2336), .ZN(n_5_2085));
   INV_X1 i_5_2518 (.A(n_73), .ZN(n_5_2086));
   INV_X1 i_5_2519 (.A(n_5_2340), .ZN(n_5_2087));
   INV_X1 i_5_2520 (.A(n_76), .ZN(n_5_2091));
   NAND2_X1 i_5_2521 (.A1(n_5_2340), .A2(n_76), .ZN(n_5_2092));
   INV_X1 i_5_2522 (.A(n_5_2344), .ZN(n_5_2093));
   INV_X1 i_5_2523 (.A(n_75), .ZN(n_5_2094));
   NAND2_X1 i_5_2524 (.A1(n_5_2093), .A2(n_5_2094), .ZN(n_5_2095));
   NAND2_X1 i_5_2525 (.A1(n_5_2344), .A2(n_75), .ZN(n_5_2096));
   INV_X1 i_5_2526 (.A(n_5_2347), .ZN(n_5_2097));
   INV_X1 i_5_2527 (.A(n_61), .ZN(n_5_2098));
   NAND2_X1 i_5_2528 (.A1(n_5_2097), .A2(n_5_2098), .ZN(n_5_2099));
   NAND2_X1 i_5_2529 (.A1(n_5_2347), .A2(n_61), .ZN(n_5_2100));
   NAND2_X1 i_5_2530 (.A1(n_5_2354), .A2(n_53), .ZN(n_5_2101));
   INV_X1 i_5_2531 (.A(n_5_2354), .ZN(n_5_2102));
   NAND2_X1 i_5_2532 (.A1(n_5_2102), .A2(n_5_2081), .ZN(n_5_2103));
   INV_X1 i_5_2533 (.A(n_5_2096), .ZN(n_5_2104));
   INV_X1 i_5_2534 (.A(n_5_2100), .ZN(n_5_2105));
   INV_X1 i_5_2535 (.A(n_5_2095), .ZN(n_5_2106));
   AOI21_X1 i_5_2536 (.A(n_5_2106), .B1(n_5_2281), .B2(n_5_2096), .ZN(n_5_2107));
   NAND2_X1 i_5_2537 (.A1(n_5_2279), .A2(n_5_2095), .ZN(n_5_2108));
   NAND3_X1 i_5_2538 (.A1(n_5_2108), .A2(n_5_2100), .A3(n_5_2096), .ZN(n_5_2109));
   INV_X1 i_5_2539 (.A(n_5_2109), .ZN(n_5_2111));
   NAND2_X1 i_5_2540 (.A1(n_5_2101), .A2(n_5_2099), .ZN(n_5_2112));
   OAI21_X1 i_5_2541 (.A(n_5_2103), .B1(n_5_2111), .B2(n_5_2112), .ZN(n_5_2113));
   XNOR2_X1 i_5_2542 (.A(n_5_2347), .B(n_61), .ZN(n_5_2114));
   XNOR2_X1 i_5_2543 (.A(n_5_2149), .B(n_5_2114), .ZN(n_5_2115));
   XNOR2_X1 i_5_2544 (.A(n_5_2354), .B(n_53), .ZN(n_5_2117));
   XNOR2_X1 i_5_2545 (.A(n_5_2594), .B(n_5_2117), .ZN(n_5_2262));
   XNOR2_X1 i_5_2546 (.A(n_53), .B(n_5_2082), .ZN(n_5_2118));
   XNOR2_X1 i_5_2547 (.A(n_5_2113), .B(n_5_2118), .ZN(n_5_2119));
   XOR2_X1 i_5_2548 (.A(n_5_2121), .B(n_5_2122), .Z(n_5_2120));
   NAND2_X1 i_5_2549 (.A1(n_5_2293), .A2(n_5_2577), .ZN(n_5_2121));
   NAND2_X1 i_5_2550 (.A1(n_5_2865), .A2(m[0]), .ZN(n_5_2122));
   XNOR2_X1 i_5_2551 (.A(n_5_2597), .B(n_5_2125), .ZN(n_5_2123));
   INV_X1 i_5_2552 (.A(n_5_2124), .ZN(n_5_2263));
   NAND3_X1 i_5_2553 (.A1(n_5_2306), .A2(n_5_2574), .A3(n_5_2126), .ZN(n_5_2124));
   NAND2_X1 i_5_2554 (.A1(n_5_2220), .A2(n_5_2306), .ZN(n_5_2264));
   NAND2_X1 i_5_2555 (.A1(n_5_2140), .A2(n_5_2131), .ZN(n_5_2265));
   NAND2_X1 i_5_2556 (.A1(n_5_2133), .A2(n_5_2132), .ZN(n_5_2125));
   NAND2_X1 i_5_2557 (.A1(n_5_2574), .A2(n_5_2126), .ZN(n_5_2266));
   NAND2_X1 i_5_2558 (.A1(n_5_2570), .A2(n_5_2866), .ZN(n_5_2126));
   XNOR2_X1 i_5_2559 (.A(n_5_2300), .B(n_5_2127), .ZN(n_5_3393));
   XNOR2_X1 i_5_2560 (.A(n_5_2896), .B(n_60), .ZN(n_5_2127));
   NAND2_X1 i_5_1611 (.A1(n_5_2194), .A2(n_5_2136), .ZN(n_5_2267));
   NOR2_X1 i_5_2562 (.A1(n_5_2318), .A2(n_5_2129), .ZN(n_5_2128));
   AOI21_X1 i_5_2563 (.A(n_5_2142), .B1(n_5_2141), .B2(n_5_2136), .ZN(n_5_2129));
   NAND2_X1 i_5_2564 (.A1(n_5_2164), .A2(n_5_2130), .ZN(n_5_4071));
   NAND2_X1 i_5_2565 (.A1(n_5_2279), .A2(n_5_2151), .ZN(n_5_2130));
   OAI21_X1 i_5_2566 (.A(n_5_2131), .B1(n_5_2802), .B2(n_5_2150), .ZN(n_5_2268));
   AND2_X1 i_5_2567 (.A1(n_5_2821), .A2(n_5_2132), .ZN(n_5_2131));
   NAND2_X1 i_5_2568 (.A1(n_5_2803), .A2(n_66), .ZN(n_5_2132));
   INV_X1 i_5_2569 (.A(n_5_2802), .ZN(n_5_2133));
   INV_X1 i_5_2570 (.A(n_5_2308), .ZN(n_5_2134));
   AOI21_X1 i_5_2571 (.A(n_5_2139), .B1(n_5_2312), .B2(n_5_2138), .ZN(n_5_2135));
   NAND2_X1 i_5_2572 (.A1(n_5_3130), .A2(n_55), .ZN(n_5_2136));
   NOR2_X1 i_5_2573 (.A1(n_5_3130), .A2(n_55), .ZN(n_5_2137));
   NAND2_X1 i_5_2574 (.A1(n_5_2087), .A2(n_5_2091), .ZN(n_5_2138));
   INV_X1 i_5_2575 (.A(n_5_2092), .ZN(n_5_2139));
   INV_X1 i_5_2576 (.A(n_5_2223), .ZN(n_5_2269));
   OAI21_X1 i_5_2577 (.A(n_5_2133), .B1(n_5_2597), .B2(n_5_2125), .ZN(n_5_2140));
   NAND3_X1 i_5_2578 (.A1(n_5_2231), .A2(n_5_2194), .A3(n_5_2244), .ZN(n_5_2141));
   XNOR2_X1 i_5_2579 (.A(n_5_2336), .B(n_73), .ZN(n_5_2142));
   XNOR2_X1 i_5_2580 (.A(n_5_2336), .B(n_73), .ZN(n_5_2143));
   NAND3_X1 i_5_2581 (.A1(n_5_2231), .A2(n_5_2194), .A3(n_5_2244), .ZN(n_5_2144));
   INV_X1 i_5_2582 (.A(n_5_3185), .ZN(n_5_2145));
   NAND2_X1 i_5_2583 (.A1(n_5_2104), .A2(n_5_2095), .ZN(n_5_2146));
   INV_X1 i_5_2584 (.A(n_5_2279), .ZN(n_5_2147));
   INV_X1 i_5_2585 (.A(n_5_2095), .ZN(n_5_2148));
   OAI21_X1 i_5_2586 (.A(n_5_2146), .B1(n_5_2147), .B2(n_5_2148), .ZN(n_5_2149));
   NAND2_X1 i_5_2587 (.A1(n_5_2812), .A2(n_5_2579), .ZN(n_5_2150));
   XNOR2_X1 i_5_2588 (.A(n_5_2344), .B(n_75), .ZN(n_5_2151));
   INV_X1 i_5_2589 (.A(n_75), .ZN(n_5_2152));
   XNOR2_X1 i_5_2590 (.A(n_5_2344), .B(n_5_2152), .ZN(n_5_2163));
   NAND3_X1 i_5_2591 (.A1(n_5_2163), .A2(n_5_2135), .A3(n_5_2991), .ZN(n_5_2164));
   NOR2_X1 i_5_2592 (.A1(n_5_2597), .A2(n_5_2125), .ZN(n_5_2171));
   NAND2_X1 i_5_2593 (.A1(n_5_2171), .A2(n_5_2823), .ZN(n_5_2172));
   XNOR2_X1 i_5_2594 (.A(n_5_2823), .B(n_5_2133), .ZN(n_5_2173));
   OAI21_X1 i_5_2595 (.A(n_5_2172), .B1(n_5_2173), .B2(n_5_2171), .ZN(n_5_2175));
   NAND2_X1 i_5_2596 (.A1(n_5_2316), .A2(n_5_2577), .ZN(n_5_2176));
   XNOR2_X1 i_5_2597 (.A(n_5_2303), .B(n_5_2176), .ZN(n_5_2177));
   NAND2_X1 i_5_2598 (.A1(n_5_2570), .A2(n_5_2866), .ZN(n_5_2183));
   INV_X1 i_5_2599 (.A(n_5_2183), .ZN(n_5_2193));
   INV_X1 i_5_2600 (.A(n_5_2137), .ZN(n_5_2194));
   NAND2_X1 i_5_2601 (.A1(n_5_2085), .A2(n_5_2086), .ZN(n_5_2195));
   INV_X1 i_5_2602 (.A(n_5_2137), .ZN(n_5_2200));
   NAND2_X1 i_5_2603 (.A1(n_5_2133), .A2(n_5_2226), .ZN(n_5_2201));
   INV_X1 i_5_2604 (.A(n_5_2201), .ZN(n_5_2270));
   NAND2_X1 i_5_2605 (.A1(n_5_2821), .A2(n_5_2132), .ZN(n_5_2205));
   INV_X1 i_5_2606 (.A(n_5_2205), .ZN(n_5_2215));
   OAI21_X1 i_5_2607 (.A(n_5_2215), .B1(n_5_2224), .B2(n_5_2802), .ZN(n_5_2220));
   XOR2_X1 i_5_2608 (.A(n_5_2809), .B(n_5_2246), .Z(n_5_2222));
   AOI21_X1 i_5_2609 (.A(n_5_2301), .B1(n_5_2315), .B2(n_5_2794), .ZN(n_5_2223));
   NAND2_X1 i_5_2610 (.A1(n_5_2596), .A2(n_5_2226), .ZN(n_5_2224));
   OR2_X1 i_5_2611 (.A1(n_5_2812), .A2(n_5_2579), .ZN(n_5_2226));
   NOR2_X1 i_5_2612 (.A1(n_5_2812), .A2(n_5_2579), .ZN(n_5_2227));
   NAND2_X1 i_5_2613 (.A1(n_5_2896), .A2(n_60), .ZN(n_5_2230));
   NAND2_X1 i_5_2614 (.A1(n_5_3255), .A2(n_5_3256), .ZN(n_5_2231));
   NAND2_X1 i_5_2615 (.A1(n_5_2083), .A2(n_5_2084), .ZN(n_5_2244));
   NAND2_X1 i_5_2616 (.A1(n_5_2083), .A2(n_5_2084), .ZN(n_5_2271));
   AOI21_X1 i_5_2617 (.A(n_5_2301), .B1(n_5_2314), .B2(n_5_2794), .ZN(n_5_2246));
   NAND2_X1 i_5_2618 (.A1(n_5_2315), .A2(n_5_2794), .ZN(n_5_2272));
   XNOR2_X1 i_5_2619 (.A(n_5_2314), .B(n_5_2792), .ZN(n_5_2273));
   INV_X1 i_5_2620 (.A(n_5_2896), .ZN(n_5_2274));
   INV_X1 i_5_2621 (.A(n_5_2193), .ZN(n_5_2275));
   NAND2_X1 i_5_2622 (.A1(n_5_2274), .A2(n_5_2275), .ZN(n_5_2276));
   INV_X1 i_5_2623 (.A(n_60), .ZN(n_5_2277));
   NAND2_X1 i_5_2624 (.A1(n_5_2275), .A2(n_5_2277), .ZN(n_5_2278));
   NAND2_X1 i_5_2625 (.A1(n_5_2991), .A2(n_5_2135), .ZN(n_5_2279));
   NAND2_X1 i_5_2626 (.A1(n_5_2135), .A2(n_5_2991), .ZN(n_5_2280));
   INV_X1 i_5_2627 (.A(n_5_2280), .ZN(n_5_2281));
   NAND2_X1 i_5_2628 (.A1(n_5_2307), .A2(n_5_2136), .ZN(n_5_2282));
   INV_X1 i_5_2629 (.A(n_5_2282), .ZN(n_5_2283));
   NAND2_X1 i_5_2630 (.A1(n_5_2141), .A2(n_5_2283), .ZN(n_5_2284));
   INV_X1 i_5_2631 (.A(n_5_2284), .ZN(n_5_2285));
   INV_X1 i_5_2632 (.A(n_76), .ZN(n_5_2286));
   XNOR2_X1 i_5_2633 (.A(n_5_2340), .B(n_5_2286), .ZN(n_5_2287));
   NAND2_X1 i_5_2634 (.A1(n_5_2285), .A2(n_5_2287), .ZN(n_5_2288));
   XNOR2_X1 i_5_2635 (.A(n_76), .B(n_5_2086), .ZN(n_5_2289));
   XNOR2_X1 i_5_2636 (.A(n_5_2340), .B(n_5_2289), .ZN(n_5_2290));
   MUX2_X1 i_5_2637 (.A(n_5_2287), .B(n_5_2290), .S(n_5_2085), .Z(n_5_2291));
   OAI21_X1 i_5_2638 (.A(n_5_2288), .B1(n_5_2291), .B2(n_5_2285), .ZN(n_5_2292));
   OR2_X1 i_5_2639 (.A1(n_5_2886), .A2(n_5_2568), .ZN(n_5_2293));
   NAND2_X1 i_5_2640 (.A1(n_5_2865), .A2(m[0]), .ZN(n_5_2294));
   INV_X1 i_5_2641 (.A(n_5_2294), .ZN(n_5_2295));
   NAND2_X1 i_5_2642 (.A1(n_5_2133), .A2(n_5_2226), .ZN(n_5_2296));
   NOR2_X1 i_5_2643 (.A1(n_5_2296), .A2(n_5_2223), .ZN(n_5_2297));
   OAI21_X1 i_5_2644 (.A(n_5_2304), .B1(n_5_2297), .B2(n_5_2268), .ZN(n_5_2298));
   INV_X1 i_5_2645 (.A(n_5_2193), .ZN(n_5_2299));
   NAND2_X1 i_5_2646 (.A1(n_5_2298), .A2(n_5_2299), .ZN(n_5_2300));
   INV_X1 i_5_2647 (.A(n_5_2793), .ZN(n_5_2301));
   NAND2_X1 i_5_2648 (.A1(n_5_2105), .A2(n_5_2099), .ZN(n_5_2302));
   XNOR2_X1 i_5_2649 (.A(n_5_2867), .B(n_5_3329), .ZN(n_5_2303));
   INV_X1 i_5_2650 (.A(n_5_2305), .ZN(n_5_2304));
   NAND2_X1 i_5_2651 (.A1(n_5_2574), .A2(n_5_2822), .ZN(n_5_2305));
   OR2_X1 i_5_2652 (.A1(n_5_2824), .A2(n_5_3185), .ZN(n_5_2306));
   NAND2_X1 i_5_2653 (.A1(n_5_2336), .A2(n_73), .ZN(n_5_2307));
   NAND2_X1 i_5_2654 (.A1(n_5_2195), .A2(n_5_2200), .ZN(n_5_2308));
   NAND2_X1 i_5_2655 (.A1(n_5_2136), .A2(n_5_2230), .ZN(n_5_2309));
   NAND3_X1 i_5_2656 (.A1(n_5_2200), .A2(n_5_2195), .A3(n_5_2309), .ZN(n_5_2310));
   NAND2_X1 i_5_2657 (.A1(n_5_2336), .A2(n_73), .ZN(n_5_2311));
   NAND2_X1 i_5_2658 (.A1(n_5_2310), .A2(n_5_2311), .ZN(n_5_2312));
   OAI21_X1 i_5_2659 (.A(n_5_2295), .B1(n_5_2886), .B2(n_5_2568), .ZN(n_5_2313));
   AOI21_X1 i_5_2660 (.A(n_5_2806), .B1(n_5_2313), .B2(n_5_2578), .ZN(n_5_2314));
   AOI21_X1 i_5_2661 (.A(n_5_2806), .B1(n_5_2316), .B2(n_5_2578), .ZN(n_5_2315));
   OAI21_X1 i_5_2662 (.A(n_5_2295), .B1(n_5_2886), .B2(n_5_2568), .ZN(n_5_2316));
   NAND3_X1 i_5_2663 (.A1(n_5_2144), .A2(n_5_2143), .A3(n_5_2136), .ZN(n_5_2317));
   INV_X1 i_5_2664 (.A(n_5_2317), .ZN(n_5_2318));
   NAND2_X1 i_5_2665 (.A1(n_64), .A2(n_5_2835), .ZN(n_5_2319));
   NAND2_X1 i_5_2666 (.A1(n_5_2605), .A2(n_5_2352), .ZN(n_5_2320));
   NAND2_X1 i_5_2667 (.A1(n_5_2391), .A2(n_5_4209), .ZN(n_5_2321));
   NAND2_X1 i_5_2668 (.A1(n_70), .A2(n_5_2835), .ZN(n_5_2322));
   NAND2_X1 i_5_2669 (.A1(n_5_2689), .A2(n_5_2352), .ZN(n_5_2323));
   NAND2_X1 i_5_2670 (.A1(n_62), .A2(n_5_2835), .ZN(n_5_2324));
   INV_X1 i_5_2671 (.A(n_5_2324), .ZN(n_5_2325));
   AOI21_X1 i_5_2672 (.A(n_5_2325), .B1(n_5_2385), .B2(n_5_4209), .ZN(n_5_2326));
   NAND2_X1 i_5_2673 (.A1(n_5_2444), .A2(n_5_4209), .ZN(n_5_2327));
   NAND2_X1 i_5_2674 (.A1(n_5_2767), .A2(n_5_2352), .ZN(n_5_2328));
   NAND2_X1 i_5_2675 (.A1(n_48), .A2(n_5_2835), .ZN(n_5_2329));
   NAND2_X1 i_5_2676 (.A1(n_74), .A2(n_5_2355), .ZN(n_5_2330));
   NAND2_X1 i_5_2677 (.A1(n_77), .A2(n_5_2355), .ZN(n_5_2331));
   INV_X1 i_5_2678 (.A(n_5_2331), .ZN(n_5_2332));
   NAND2_X1 i_5_2679 (.A1(n_5_2671), .A2(n_5_2352), .ZN(n_5_2333));
   NAND2_X1 i_5_2680 (.A1(n_49), .A2(n_5_2355), .ZN(n_5_2334));
   INV_X1 i_5_2681 (.A(n_5_2334), .ZN(n_5_2335));
   NAND2_X1 i_5_2682 (.A1(n_5_2333), .A2(n_5_4181), .ZN(n_5_2336));
   NAND2_X1 i_5_2683 (.A1(n_5_2484), .A2(n_5_4209), .ZN(n_5_2337));
   NAND2_X1 i_5_2684 (.A1(n_5_2610), .A2(n_5_2352), .ZN(n_5_2338));
   NAND2_X1 i_5_2685 (.A1(n_5_4200), .A2(n_5_2355), .ZN(n_5_2339));
   NAND3_X1 i_5_2686 (.A1(n_5_2337), .A2(n_5_2338), .A3(n_5_2339), .ZN(n_5_2340));
   NAND2_X1 i_5_2687 (.A1(n_5_2612), .A2(n_5_2352), .ZN(n_5_2341));
   NAND2_X1 i_5_2688 (.A1(n_5_2364), .A2(n_5_4209), .ZN(n_5_2342));
   NAND2_X1 i_5_2689 (.A1(n_51), .A2(n_5_2355), .ZN(n_5_2343));
   NAND3_X1 i_5_2690 (.A1(n_5_2341), .A2(n_5_2342), .A3(n_5_2343), .ZN(n_5_2344));
   NAND2_X1 i_5_2691 (.A1(n_5_2615), .A2(n_5_2352), .ZN(n_5_2345));
   NAND2_X1 i_5_2692 (.A1(n_5_2366), .A2(n_5_4209), .ZN(n_5_2346));
   NAND3_X1 i_5_2693 (.A1(n_5_2345), .A2(n_5_2346), .A3(n_5_2350), .ZN(n_5_2347));
   INV_X1 i_5_2694 (.A(r[0]), .ZN(n_5_2348));
   NAND2_X1 i_5_2695 (.A1(r[1]), .A2(n_5_2348), .ZN(n_5_4072));
   NAND2_X1 i_5_2696 (.A1(n_5_2368), .A2(n_5_4209), .ZN(n_5_2349));
   NAND2_X1 i_5_2697 (.A1(n_52), .A2(n_5_2355), .ZN(n_5_2350));
   INV_X1 i_5_2698 (.A(n_5_2350), .ZN(n_5_2351));
   NOR2_X1 i_5_2699 (.A1(r[1]), .A2(n_5_2348), .ZN(n_5_2352));
   AOI21_X1 i_5_2700 (.A(n_5_2351), .B1(n_5_2619), .B2(n_5_2352), .ZN(n_5_2353));
   NAND2_X1 i_5_2701 (.A1(n_5_2349), .A2(n_5_2353), .ZN(n_5_2354));
   BUF_X1 rt_shieldBuf__2__2__2 (.A(n_5_2835), .Z(n_5_2355));
   XNOR2_X1 i_5_2702 (.A(r[1]), .B(r[0]), .ZN(n_5_2356));
   XNOR2_X1 i_5_2703 (.A(r[1]), .B(r[0]), .ZN(n_5_2357));
   NAND2_X1 i_5_2704 (.A1(n_5_2835), .A2(n_67), .ZN(n_5_2358));
   INV_X1 i_5_2705 (.A(n_5_4072), .ZN(n_5_2359));
   NAND2_X1 i_5_2706 (.A1(n_5_2357), .A2(n_71), .ZN(n_5_2360));
   XNOR2_X1 i_5_2707 (.A(n_5_2381), .B(n_5_2362), .ZN(n_5_2361));
   OAI21_X1 i_5_2708 (.A(n_5_2384), .B1(n_56), .B2(n_63), .ZN(n_5_2362));
   NOR2_X1 i_5_2709 (.A1(n_5_2424), .A2(n_5_2398), .ZN(n_5_2363));
   AOI21_X1 i_5_2710 (.A(n_5_2370), .B1(n_5_2376), .B2(n_5_2365), .ZN(n_5_2364));
   OAI21_X1 i_5_2711 (.A(n_5_2452), .B1(n_75), .B2(n_5_4200), .ZN(n_5_2365));
   XNOR2_X1 i_5_2712 (.A(n_5_2370), .B(n_5_2367), .ZN(n_5_2366));
   OAI22_X1 i_5_2713 (.A1(n_53), .A2(n_52), .B1(n_5_2377), .B2(n_5_2374), 
      .ZN(n_5_2367));
   XNOR2_X1 i_5_2714 (.A(n_54), .B(n_5_2369), .ZN(n_5_2368));
   OAI222_X1 i_5_2715 (.A1(n_53), .A2(n_5_2371), .B1(n_5_2377), .B2(n_5_2374), 
      .C1(n_52), .C2(n_5_2370), .ZN(n_5_2369));
   INV_X1 i_5_2716 (.A(n_5_2371), .ZN(n_5_2370));
   OAI211_X1 i_5_2717 (.A(n_61), .B(n_5_2452), .C1(n_75), .C2(n_5_4200), 
      .ZN(n_5_2371));
   INV_X1 i_5_2718 (.A(n_5_2373), .ZN(n_5_2372));
   NAND2_X1 i_5_2719 (.A1(n_73), .A2(n_77), .ZN(n_5_2373));
   INV_X1 i_5_2720 (.A(n_52), .ZN(n_5_2374));
   INV_X1 i_5_2721 (.A(n_75), .ZN(n_5_2375));
   INV_X1 i_5_2722 (.A(n_61), .ZN(n_5_2376));
   INV_X1 i_5_2723 (.A(n_53), .ZN(n_5_2377));
   NAND2_X1 i_5_2724 (.A1(n_5_2400), .A2(n_5_2587), .ZN(n_5_2378));
   INV_X1 i_5_2725 (.A(n_5_2460), .ZN(n_5_2379));
   NOR2_X1 i_5_2726 (.A1(n_62), .A2(n_69), .ZN(n_5_2380));
   INV_X1 i_5_2727 (.A(n_5_2495), .ZN(n_5_2381));
   INV_X1 i_5_2728 (.A(n_5_4441), .ZN(n_5_2382));
   INV_X1 i_5_2729 (.A(n_55), .ZN(n_5_2383));
   NAND2_X1 i_5_2730 (.A1(n_63), .A2(n_56), .ZN(n_5_2384));
   NAND2_X1 i_5_2731 (.A1(n_5_2506), .A2(n_5_2386), .ZN(n_5_2385));
   NAND3_X1 i_5_2732 (.A1(n_5_2490), .A2(n_5_2502), .A3(n_5_2489), .ZN(n_5_2386));
   INV_X1 i_5_2733 (.A(n_64), .ZN(n_5_2387));
   INV_X1 i_5_2734 (.A(n_66), .ZN(n_5_2388));
   INV_X1 i_5_2735 (.A(n_5_2379), .ZN(n_5_2389));
   INV_X1 i_5_2736 (.A(n_5_2380), .ZN(n_5_2390));
   NAND2_X1 i_5_2737 (.A1(n_5_3838), .A2(n_5_2537), .ZN(n_5_4073));
   NAND2_X1 i_5_2738 (.A1(n_5_2392), .A2(n_5_2394), .ZN(n_5_2391));
   NAND3_X1 i_5_2739 (.A1(n_5_2485), .A2(n_5_2393), .A3(n_5_2580), .ZN(n_5_2392));
   NAND2_X1 i_5_2740 (.A1(n_5_2502), .A2(n_5_2543), .ZN(n_5_2393));
   NAND2_X1 i_5_2741 (.A1(n_5_2508), .A2(n_5_2395), .ZN(n_5_2394));
   NAND3_X1 i_5_2742 (.A1(n_5_2497), .A2(n_5_2580), .A3(n_5_2522), .ZN(n_5_2395));
   INV_X1 i_5_2743 (.A(n_59), .ZN(n_5_2396));
   NAND3_X1 i_5_2744 (.A1(n_5_2580), .A2(n_66), .A3(n_64), .ZN(n_5_2397));
   INV_X1 i_5_2745 (.A(n_5_2422), .ZN(n_5_2398));
   NAND2_X1 i_5_2746 (.A1(n_5_2449), .A2(n_5_2401), .ZN(n_5_2399));
   NAND2_X1 i_5_2747 (.A1(n_5_4444), .A2(n_5_2401), .ZN(n_5_2400));
   INV_X1 i_5_2748 (.A(n_5_2402), .ZN(n_5_2401));
   NOR2_X1 i_5_2749 (.A1(n_74), .A2(n_55), .ZN(n_5_2402));
   NAND2_X1 i_5_2750 (.A1(n_5_2404), .A2(n_5_2419), .ZN(n_5_2403));
   INV_X1 i_5_2751 (.A(n_5_2372), .ZN(n_5_2404));
   INV_X1 i_5_2752 (.A(n_5_2413), .ZN(n_5_2405));
   NAND2_X1 i_5_2753 (.A1(n_5_2407), .A2(n_5_2408), .ZN(n_5_2406));
   INV_X1 i_5_2754 (.A(n_5_2441), .ZN(n_5_2407));
   INV_X1 i_5_2755 (.A(n_5_2375), .ZN(n_5_2408));
   INV_X1 i_5_2756 (.A(n_50), .ZN(n_5_2409));
   INV_X1 i_5_2757 (.A(n_75), .ZN(n_5_2410));
   OAI21_X1 i_5_2758 (.A(n_5_2440), .B1(n_5_2425), .B2(n_5_2426), .ZN(n_5_2411));
   NAND3_X1 i_5_2759 (.A1(n_5_2422), .A2(n_5_2373), .A3(n_5_2413), .ZN(n_5_2412));
   NAND3_X1 i_5_2760 (.A1(n_5_2449), .A2(n_5_2841), .A3(n_5_2419), .ZN(n_5_2413));
   NOR2_X1 i_5_2761 (.A1(n_62), .A2(n_69), .ZN(n_5_2414));
   NOR2_X1 i_5_2762 (.A1(n_48), .A2(n_60), .ZN(n_5_2415));
   NAND2_X1 i_5_2763 (.A1(n_5_2529), .A2(n_5_2540), .ZN(n_5_2416));
   INV_X1 i_5_2764 (.A(n_67), .ZN(n_5_2417));
   INV_X1 i_5_2765 (.A(n_58), .ZN(n_5_2418));
   NAND2_X1 i_5_2766 (.A1(n_5_2420), .A2(n_5_2421), .ZN(n_5_2419));
   INV_X1 i_5_2767 (.A(n_77), .ZN(n_5_2420));
   INV_X1 i_5_2768 (.A(n_73), .ZN(n_5_2421));
   NAND2_X1 i_5_2769 (.A1(n_49), .A2(n_76), .ZN(n_5_2422));
   INV_X1 i_5_2770 (.A(n_5_2424), .ZN(n_5_2423));
   NOR2_X1 i_5_2771 (.A1(n_49), .A2(n_76), .ZN(n_5_2424));
   NOR2_X1 i_5_2772 (.A1(n_5_2441), .A2(n_5_2375), .ZN(n_5_2425));
   NOR2_X1 i_5_2773 (.A1(n_50), .A2(n_75), .ZN(n_5_2426));
   INV_X1 i_5_2774 (.A(n_62), .ZN(n_5_2427));
   INV_X1 i_5_2775 (.A(n_5_2474), .ZN(n_5_2428));
   INV_X1 i_5_2776 (.A(n_5_2396), .ZN(n_5_2429));
   NAND2_X1 i_5_2777 (.A1(n_5_2428), .A2(n_5_2429), .ZN(n_5_2430));
   INV_X1 i_5_2778 (.A(n_5_3834), .ZN(n_5_2431));
   INV_X1 i_5_2779 (.A(n_5_3835), .ZN(n_5_2432));
   NAND2_X1 i_5_2780 (.A1(n_5_2431), .A2(n_5_2432), .ZN(n_5_2433));
   NAND2_X1 i_5_2781 (.A1(n_71), .A2(n_65), .ZN(n_5_2434));
   NAND2_X1 i_5_2782 (.A1(n_72), .A2(n_59), .ZN(n_5_2435));
   INV_X1 i_5_2783 (.A(n_5_3835), .ZN(n_5_2436));
   NAND2_X1 i_5_2784 (.A1(n_5_2550), .A2(n_5_2436), .ZN(n_5_2437));
   INV_X1 i_5_2785 (.A(n_5_2399), .ZN(n_5_2438));
   NAND2_X1 i_5_2786 (.A1(n_5_2387), .A2(n_5_2388), .ZN(n_5_2439));
   NAND2_X1 i_5_2787 (.A1(n_5_2412), .A2(n_5_2423), .ZN(n_5_2440));
   INV_X1 i_5_2788 (.A(n_50), .ZN(n_5_2441));
   INV_X1 i_5_2789 (.A(n_5_2375), .ZN(n_5_2442));
   NOR2_X1 i_5_2790 (.A1(n_5_2382), .A2(n_5_2415), .ZN(n_5_2443));
   XNOR2_X1 i_5_2791 (.A(n_5_2876), .B(n_5_2443), .ZN(n_5_2444));
   NAND2_X1 i_5_2792 (.A1(n_5_2399), .A2(n_5_2403), .ZN(n_5_2445));
   NAND2_X1 i_5_2793 (.A1(n_48), .A2(n_60), .ZN(n_5_2446));
   INV_X1 i_5_2794 (.A(n_5_2446), .ZN(n_5_2447));
   AOI21_X1 i_5_2795 (.A(n_5_2447), .B1(n_74), .B2(n_55), .ZN(n_5_2448));
   NAND2_X1 i_5_2796 (.A1(n_5_2519), .A2(n_5_2448), .ZN(n_5_2449));
   NAND2_X1 i_5_2797 (.A1(n_5_2423), .A2(n_5_2412), .ZN(n_5_2450));
   NAND2_X1 i_5_2798 (.A1(n_50), .A2(n_5_2442), .ZN(n_5_2451));
   NAND2_X1 i_5_2799 (.A1(n_5_2450), .A2(n_5_2451), .ZN(n_5_2452));
   NAND2_X1 i_5_2800 (.A1(n_72), .A2(n_59), .ZN(n_5_2453));
   INV_X1 i_5_2801 (.A(n_5_2396), .ZN(n_5_2454));
   NAND2_X1 i_5_2802 (.A1(n_67), .A2(n_58), .ZN(n_5_2455));
   INV_X1 i_5_2803 (.A(n_5_2417), .ZN(n_5_2456));
   INV_X1 i_5_2804 (.A(n_5_2418), .ZN(n_5_2457));
   OAI21_X1 i_5_2805 (.A(n_5_2455), .B1(n_5_2456), .B2(n_5_2457), .ZN(n_5_2458));
   OAI21_X1 i_5_2806 (.A(n_5_2439), .B1(n_70), .B2(n_68), .ZN(n_5_2459));
   NAND2_X1 i_5_2807 (.A1(n_62), .A2(n_69), .ZN(n_5_2460));
   INV_X1 i_5_2808 (.A(n_5_2427), .ZN(n_5_2461));
   NAND2_X1 i_5_2809 (.A1(n_70), .A2(n_5_2546), .ZN(n_5_2462));
   INV_X1 i_5_2810 (.A(n_68), .ZN(n_5_2463));
   NOR2_X1 i_5_2811 (.A1(n_5_2427), .A2(n_5_2463), .ZN(n_5_2464));
   NAND2_X1 i_5_2812 (.A1(n_70), .A2(n_5_2464), .ZN(n_5_2465));
   NAND2_X1 i_5_2813 (.A1(n_69), .A2(n_62), .ZN(n_5_2466));
   NAND3_X1 i_5_2814 (.A1(n_5_2462), .A2(n_5_2465), .A3(n_5_2466), .ZN(n_5_2467));
   INV_X1 i_5_2815 (.A(n_5_2467), .ZN(n_5_2468));
   NAND2_X1 i_5_2816 (.A1(n_5_2434), .A2(n_5_2430), .ZN(n_5_2469));
   NAND3_X1 i_5_2817 (.A1(n_5_2435), .A2(n_5_2536), .A3(n_5_2437), .ZN(n_5_2470));
   NAND2_X1 i_5_2818 (.A1(n_5_2474), .A2(n_5_2396), .ZN(n_5_2471));
   NAND3_X1 i_5_2819 (.A1(n_5_2536), .A2(n_5_2437), .A3(n_5_2435), .ZN(n_5_2472));
   NAND2_X1 i_5_2820 (.A1(n_5_2474), .A2(n_5_2396), .ZN(n_5_2473));
   INV_X1 i_5_2821 (.A(n_72), .ZN(n_5_2474));
   NAND2_X1 i_5_2822 (.A1(n_5_2472), .A2(n_5_2473), .ZN(n_5_2475));
   INV_X1 i_5_2823 (.A(n_5_2472), .ZN(n_5_2476));
   INV_X1 i_5_2824 (.A(n_65), .ZN(n_5_2477));
   NAND2_X1 i_5_2825 (.A1(n_5_2476), .A2(n_5_2482), .ZN(n_5_2478));
   OAI21_X1 i_5_2826 (.A(n_5_2478), .B1(n_5_2481), .B2(n_5_2476), .ZN(n_5_2479));
   XNOR2_X1 i_5_2827 (.A(n_71), .B(n_5_2477), .ZN(n_5_2480));
   XNOR2_X1 i_5_2828 (.A(n_5_2480), .B(n_5_2473), .ZN(n_5_2481));
   XNOR2_X1 i_5_2829 (.A(n_71), .B(n_5_2477), .ZN(n_5_2482));
   NAND2_X1 i_5_2830 (.A1(n_5_2819), .A2(n_5_2411), .ZN(n_5_2483));
   INV_X1 i_5_2831 (.A(n_5_2483), .ZN(n_5_2484));
   NAND3_X1 i_5_2832 (.A1(n_5_2539), .A2(n_5_2540), .A3(n_5_2538), .ZN(n_5_2485));
   NAND2_X1 i_5_2833 (.A1(n_5_2417), .A2(n_5_2418), .ZN(n_5_2486));
   NAND2_X1 i_5_2834 (.A1(n_5_2902), .A2(n_5_2527), .ZN(n_5_2487));
   INV_X1 i_5_2835 (.A(n_5_2901), .ZN(n_5_2488));
   NAND2_X1 i_5_2836 (.A1(n_5_2503), .A2(n_5_2543), .ZN(n_5_2489));
   NAND2_X1 i_5_2837 (.A1(n_5_2389), .A2(n_5_2390), .ZN(n_5_2490));
   INV_X1 i_5_2838 (.A(n_70), .ZN(n_5_2491));
   INV_X1 i_5_2839 (.A(n_68), .ZN(n_5_2492));
   NAND4_X1 i_5_2840 (.A1(n_5_2491), .A2(n_5_2389), .A3(n_5_2390), .A4(n_5_2492), 
      .ZN(n_5_2493));
   NAND3_X1 i_5_2841 (.A1(n_5_2543), .A2(n_5_2389), .A3(n_5_2390), .ZN(n_5_2494));
   NAND2_X1 i_5_2842 (.A1(n_57), .A2(m[0]), .ZN(n_5_2495));
   INV_X1 i_5_2843 (.A(n_5_2424), .ZN(n_5_4074));
   NAND2_X1 i_5_2844 (.A1(n_5_2409), .A2(n_5_2410), .ZN(n_5_2496));
   NAND3_X1 i_5_2845 (.A1(n_5_2529), .A2(n_5_2499), .A3(n_5_2500), .ZN(n_5_2497));
   NAND2_X1 i_5_2846 (.A1(n_5_2417), .A2(n_5_2418), .ZN(n_5_2498));
   NAND3_X1 i_5_2847 (.A1(n_5_2470), .A2(n_5_2523), .A3(n_5_2471), .ZN(n_5_2499));
   NAND2_X1 i_5_2848 (.A1(n_71), .A2(n_65), .ZN(n_5_2500));
   OR2_X1 i_5_2849 (.A1(n_70), .A2(n_68), .ZN(n_5_2501));
   OR2_X1 i_5_2850 (.A1(n_70), .A2(n_68), .ZN(n_5_2502));
   NAND2_X1 i_5_2851 (.A1(n_5_2554), .A2(n_5_2580), .ZN(n_5_2503));
   NAND3_X1 i_5_2852 (.A1(n_5_2554), .A2(n_5_2493), .A3(n_5_2580), .ZN(n_5_2504));
   NAND2_X1 i_5_2853 (.A1(n_5_2494), .A2(n_5_2493), .ZN(n_5_2505));
   NAND2_X1 i_5_2854 (.A1(n_5_2504), .A2(n_5_2505), .ZN(n_5_2506));
   NAND2_X1 i_5_2855 (.A1(n_5_2433), .A2(n_5_2495), .ZN(n_5_2507));
   INV_X1 i_5_2856 (.A(n_5_2544), .ZN(n_5_2508));
   NAND3_X1 i_5_2857 (.A1(n_5_2523), .A2(n_5_2470), .A3(n_5_2471), .ZN(n_5_2509));
   NAND2_X1 i_5_2858 (.A1(n_71), .A2(n_65), .ZN(n_5_2510));
   INV_X1 i_5_2859 (.A(n_5_2510), .ZN(n_5_2511));
   AOI21_X1 i_5_2860 (.A(n_5_2511), .B1(n_67), .B2(n_58), .ZN(n_5_2512));
   NAND2_X1 i_5_2861 (.A1(n_5_2509), .A2(n_5_2512), .ZN(n_5_2513));
   NAND3_X1 i_5_2862 (.A1(n_5_2826), .A2(n_5_2828), .A3(n_5_2827), .ZN(n_5_4075));
   NOR2_X1 i_5_2863 (.A1(n_5_2414), .A2(n_5_2415), .ZN(n_5_4076));
   NAND3_X1 i_5_2864 (.A1(n_5_2459), .A2(n_5_2543), .A3(n_5_2460), .ZN(n_5_4077));
   NAND3_X1 i_5_2865 (.A1(n_5_2827), .A2(n_5_2826), .A3(n_5_2828), .ZN(n_5_2514));
   NAND3_X1 i_5_2866 (.A1(n_5_2543), .A2(n_5_2459), .A3(n_5_2460), .ZN(n_5_2515));
   INV_X1 i_5_2867 (.A(n_5_2414), .ZN(n_5_2516));
   NAND2_X1 i_5_2868 (.A1(n_5_2515), .A2(n_5_2516), .ZN(n_5_2517));
   NOR2_X1 i_5_2869 (.A1(n_5_2517), .A2(n_5_2415), .ZN(n_5_2518));
   NAND2_X1 i_5_2870 (.A1(n_5_2514), .A2(n_5_2518), .ZN(n_5_2519));
   NAND2_X1 i_5_2871 (.A1(n_5_2535), .A2(n_5_2439), .ZN(n_5_2520));
   NAND2_X1 i_5_2872 (.A1(n_5_4444), .A2(n_5_2817), .ZN(n_5_2521));
   NAND2_X1 i_5_2873 (.A1(n_5_2417), .A2(n_5_2418), .ZN(n_5_2522));
   INV_X1 i_5_2874 (.A(n_5_2901), .ZN(n_5_2523));
   NAND2_X1 i_5_2875 (.A1(n_5_2475), .A2(n_5_2434), .ZN(n_5_2524));
   AOI21_X1 i_5_2876 (.A(n_5_2901), .B1(n_5_2417), .B2(n_5_2418), .ZN(n_5_2525));
   NAND2_X1 i_5_2877 (.A1(n_5_2434), .A2(n_5_2430), .ZN(n_5_2526));
   INV_X1 i_5_2878 (.A(n_5_2526), .ZN(n_5_2527));
   INV_X1 i_5_2879 (.A(n_56), .ZN(n_5_2528));
   NAND2_X1 i_5_2880 (.A1(n_67), .A2(n_58), .ZN(n_5_2529));
   NAND2_X1 i_5_2881 (.A1(n_67), .A2(n_58), .ZN(n_5_2530));
   INV_X1 i_5_2882 (.A(n_5_2530), .ZN(n_5_2531));
   OAI21_X1 i_5_2883 (.A(n_5_2461), .B1(n_70), .B2(n_68), .ZN(n_5_2532));
   NAND2_X1 i_5_2884 (.A1(n_70), .A2(n_69), .ZN(n_5_2533));
   NAND2_X1 i_5_2885 (.A1(n_68), .A2(n_69), .ZN(n_5_2534));
   NAND3_X1 i_5_2886 (.A1(n_5_2532), .A2(n_5_2533), .A3(n_5_2534), .ZN(n_5_2535));
   NAND3_X1 i_5_2887 (.A1(n_5_2548), .A2(m[0]), .A3(n_57), .ZN(n_5_2536));
   NAND2_X1 i_5_2888 (.A1(n_5_3834), .A2(n_5_2528), .ZN(n_5_2537));
   NAND3_X1 i_5_2889 (.A1(n_5_2486), .A2(n_5_2487), .A3(n_5_2488), .ZN(n_5_2538));
   NAND2_X1 i_5_2890 (.A1(n_5_2531), .A2(n_5_2522), .ZN(n_5_2539));
   NAND2_X1 i_5_2891 (.A1(n_64), .A2(n_66), .ZN(n_5_2540));
   NAND2_X1 i_5_2892 (.A1(n_64), .A2(n_66), .ZN(n_5_2541));
   NAND2_X1 i_5_2893 (.A1(n_70), .A2(n_68), .ZN(n_5_2542));
   NAND2_X1 i_5_2894 (.A1(n_70), .A2(n_68), .ZN(n_5_2543));
   NAND3_X1 i_5_2895 (.A1(n_5_2542), .A2(n_5_2501), .A3(n_5_2397), .ZN(n_5_2544));
   NAND2_X1 i_5_2896 (.A1(n_68), .A2(n_69), .ZN(n_5_2545));
   INV_X1 i_5_2897 (.A(n_5_2545), .ZN(n_5_2546));
   INV_X1 i_5_2898 (.A(n_63), .ZN(n_5_2547));
   NAND2_X1 i_5_2899 (.A1(n_5_2547), .A2(n_5_2528), .ZN(n_5_2548));
   AOI22_X1 i_5_2900 (.A1(n_5_3835), .A2(n_5_3834), .B1(n_5_2474), .B2(n_5_2396), 
      .ZN(n_5_2549));
   INV_X1 i_5_2901 (.A(n_5_3834), .ZN(n_5_2550));
   NAND3_X1 i_5_2902 (.A1(n_5_2487), .A2(n_5_2488), .A3(n_5_2486), .ZN(n_5_2551));
   INV_X1 i_5_2903 (.A(n_5_2541), .ZN(n_5_2552));
   AOI21_X1 i_5_2904 (.A(n_5_2552), .B1(n_5_2531), .B2(n_5_2522), .ZN(n_5_2553));
   NAND2_X1 i_5_2905 (.A1(n_5_2551), .A2(n_5_2553), .ZN(n_5_2554));
   INV_X1 i_5_2906 (.A(n_73), .ZN(n_5_2555));
   INV_X1 i_5_2907 (.A(n_77), .ZN(n_5_2556));
   NAND2_X1 i_5_2908 (.A1(n_5_2555), .A2(n_5_2556), .ZN(n_5_2557));
   OAI21_X1 i_5_2909 (.A(n_5_2557), .B1(n_5_2378), .B2(n_5_2372), .ZN(n_5_2558));
   NAND2_X1 i_5_2910 (.A1(n_5_4209), .A2(n_5_3329), .ZN(n_5_2559));
   INV_X1 i_5_2911 (.A(n_5_2559), .ZN(n_5_2560));
   NAND2_X1 i_5_2912 (.A1(n_5_2479), .A2(n_5_2560), .ZN(n_5_2561));
   NAND2_X1 i_5_2913 (.A1(n_5_2352), .A2(n_5_3329), .ZN(n_5_2562));
   INV_X1 i_5_2914 (.A(n_5_2562), .ZN(n_5_2563));
   NAND2_X1 i_5_2915 (.A1(n_5_2775), .A2(n_5_2563), .ZN(n_5_2564));
   INV_X1 i_5_2916 (.A(n_5_2360), .ZN(n_5_2565));
   NAND2_X1 i_5_2917 (.A1(n_5_2565), .A2(n_5_3329), .ZN(n_5_2566));
   NAND3_X1 i_5_2918 (.A1(n_5_2561), .A2(n_5_2564), .A3(n_5_2566), .ZN(n_5_2567));
   BUF_X1 rt_shieldBuf__2__2__4 (.A(n_56), .Z(n_5_2568));
   BUF_X1 rt_shieldBuf__2__2__5 (.A(n_65), .Z(n_5_2569));
   NAND3_X1 i_5_2919 (.A1(n_5_2327), .A2(n_5_2328), .A3(n_5_2329), .ZN(n_5_2570));
   INV_X1 i_5_2920 (.A(n_5_2866), .ZN(n_5_2571));
   NAND2_X1 i_5_2921 (.A1(n_5_2329), .A2(n_5_2571), .ZN(n_5_2572));
   INV_X1 i_5_2922 (.A(n_5_2572), .ZN(n_5_2573));
   NAND3_X1 i_5_2923 (.A1(n_5_2327), .A2(n_5_2328), .A3(n_5_2573), .ZN(n_5_2574));
   NAND2_X1 i_5_2924 (.A1(n_5_2586), .A2(n_5_4209), .ZN(n_5_2575));
   NAND2_X1 i_5_2925 (.A1(n_5_2738), .A2(n_5_2352), .ZN(n_5_2576));
   NAND2_X1 i_5_2926 (.A1(n_5_2886), .A2(n_5_2568), .ZN(n_5_2577));
   AOI21_X1 i_5_2927 (.A(n_5_2567), .B1(n_5_2886), .B2(n_5_2568), .ZN(n_5_2578));
   BUF_X1 rt_shieldBuf__2__2__6 (.A(n_58), .Z(n_5_2579));
   NAND2_X1 i_5_2928 (.A1(n_5_2387), .A2(n_5_2388), .ZN(n_5_2580));
   INV_X1 i_5_2929 (.A(n_5_2513), .ZN(n_5_2581));
   NAND2_X1 i_5_2930 (.A1(n_5_2387), .A2(n_5_2388), .ZN(n_5_2582));
   NAND2_X1 i_5_2931 (.A1(n_5_2582), .A2(n_5_2540), .ZN(n_5_2583));
   INV_X1 i_5_2932 (.A(n_5_2498), .ZN(n_5_2584));
   XNOR2_X1 i_5_2933 (.A(n_5_2583), .B(n_5_2584), .ZN(n_5_2585));
   OAI22_X1 i_5_2934 (.A1(n_5_2581), .A2(n_5_2585), .B1(n_5_2513), .B2(n_5_2583), 
      .ZN(n_5_2586));
   NAND2_X1 i_5_2935 (.A1(n_74), .A2(n_55), .ZN(n_5_2587));
   NAND2_X1 i_5_2936 (.A1(n_74), .A2(n_55), .ZN(n_5_2588));
   INV_X1 i_5_2937 (.A(n_5_2839), .ZN(n_5_2589));
   INV_X1 i_5_2938 (.A(n_5_2383), .ZN(n_5_2590));
   OAI21_X1 i_5_2939 (.A(n_5_2588), .B1(n_5_2589), .B2(n_5_2590), .ZN(n_5_2591));
   NAND3_X1 i_5_2940 (.A1(n_5_2591), .A2(n_5_4440), .A3(n_5_4441), .ZN(n_5_2592));
   NAND2_X1 i_5_2941 (.A1(n_5_2107), .A2(n_5_2099), .ZN(n_5_2593));
   NAND2_X1 i_5_2942 (.A1(n_5_2593), .A2(n_5_2302), .ZN(n_5_2594));
   AOI21_X1 i_5_2943 (.A(n_5_2301), .B1(n_5_2812), .B2(n_5_2579), .ZN(n_5_2595));
   NAND2_X1 i_5_2944 (.A1(n_5_2272), .A2(n_5_2595), .ZN(n_5_2596));
   AOI21_X1 i_5_2945 (.A(n_5_2227), .B1(n_5_2272), .B2(n_5_2598), .ZN(n_5_2597));
   AOI21_X1 i_5_2946 (.A(n_5_2301), .B1(n_5_2812), .B2(n_5_2579), .ZN(n_5_2598));
   BUF_X1 rt_shieldBuf__2__2__7 (.A(n_68), .Z(n_5_3185));
   XNOR2_X1 i_5_2947 (.A(n_5_2601), .B(n_5_2600), .ZN(n_5_2599));
   OAI21_X1 i_5_2948 (.A(n_5_2604), .B1(m[1]), .B2(n_63), .ZN(n_5_2600));
   INV_X1 i_5_2949 (.A(n_5_2603), .ZN(n_5_2601));
   XNOR2_X1 i_5_2950 (.A(n_5_2743), .B(n_5_2850), .ZN(n_5_2602));
   NAND2_X1 i_5_2951 (.A1(n_57), .A2(m[0]), .ZN(n_5_2603));
   NAND2_X1 i_5_2952 (.A1(n_63), .A2(m[1]), .ZN(n_5_2604));
   XNOR2_X1 i_5_2953 (.A(n_5_2685), .B(n_5_2606), .ZN(n_5_2605));
   NAND2_X1 i_5_2954 (.A1(n_5_2682), .A2(n_5_2649), .ZN(n_5_2606));
   NAND2_X1 i_5_2955 (.A1(n_5_2659), .A2(n_5_2609), .ZN(n_5_2607));
   INV_X1 i_5_2956 (.A(n_5_2784), .ZN(n_5_2608));
   NAND2_X1 i_5_2957 (.A1(n_62), .A2(m[7]), .ZN(n_5_2609));
   XNOR2_X1 i_5_2958 (.A(n_5_2633), .B(n_5_2611), .ZN(n_5_2610));
   NAND2_X1 i_5_2959 (.A1(n_5_2646), .A2(n_5_2645), .ZN(n_5_2611));
   XNOR2_X1 i_5_2960 (.A(n_5_2613), .B(n_5_2614), .ZN(n_5_2612));
   NAND2_X1 i_5_2961 (.A1(n_5_2693), .A2(n_5_2631), .ZN(n_5_2613));
   INV_X1 i_5_2962 (.A(n_5_2632), .ZN(n_5_2614));
   NAND2_X1 i_5_2963 (.A1(n_5_2618), .A2(n_5_2616), .ZN(n_5_2615));
   NAND3_X1 i_5_2964 (.A1(n_5_2617), .A2(n_5_2630), .A3(n_5_2693), .ZN(n_5_2616));
   NAND2_X1 i_5_2965 (.A1(n_5_2626), .A2(n_5_2628), .ZN(n_5_2617));
   OAI211_X1 i_5_2966 (.A(n_5_2628), .B(n_5_2626), .C1(n_5_2629), .C2(n_5_2690), 
      .ZN(n_5_2618));
   NAND2_X1 i_5_2967 (.A1(n_5_2620), .A2(n_5_2622), .ZN(n_5_2619));
   NAND2_X1 i_5_2968 (.A1(n_5_2621), .A2(n_5_2624), .ZN(n_5_2620));
   OAI21_X1 i_5_2969 (.A(n_5_2626), .B1(n_5_2629), .B2(n_5_2627), .ZN(n_5_2621));
   OAI211_X1 i_5_2970 (.A(n_5_2626), .B(n_5_2623), .C1(n_5_2663), .C2(n_5_2627), 
      .ZN(n_5_2622));
   INV_X1 i_5_2971 (.A(n_5_2624), .ZN(n_5_2623));
   XNOR2_X1 i_5_2972 (.A(m[14]), .B(n_5_2625), .ZN(n_5_2624));
   INV_X1 i_5_2973 (.A(m[15]), .ZN(n_5_2625));
   OR2_X1 i_5_2974 (.A1(n_52), .A2(m[14]), .ZN(n_5_2626));
   OAI21_X1 i_5_2975 (.A(n_5_2628), .B1(n_51), .B2(m[13]), .ZN(n_5_2627));
   NAND2_X1 i_5_2976 (.A1(n_52), .A2(m[14]), .ZN(n_5_2628));
   INV_X1 i_5_2977 (.A(n_5_2630), .ZN(n_5_2629));
   NAND2_X1 i_5_2978 (.A1(n_5_2632), .A2(n_5_2631), .ZN(n_5_2630));
   NAND2_X1 i_5_2979 (.A1(n_51), .A2(m[13]), .ZN(n_5_2631));
   OAI21_X1 i_5_2980 (.A(n_5_2646), .B1(n_5_2633), .B2(n_5_2644), .ZN(n_5_2632));
   NAND4_X1 i_5_2981 (.A1(n_5_2638), .A2(n_5_2635), .A3(n_5_2634), .A4(n_5_2723), 
      .ZN(n_5_2633));
   OAI21_X1 i_5_2982 (.A(n_5_2651), .B1(n_49), .B2(m[11]), .ZN(n_5_2634));
   OAI211_X1 i_5_2983 (.A(n_5_2642), .B(n_5_2636), .C1(n_49), .C2(m[11]), 
      .ZN(n_5_2635));
   NAND2_X1 i_5_2984 (.A1(n_5_2703), .A2(n_5_2637), .ZN(n_5_2636));
   NAND2_X1 i_5_2985 (.A1(n_48), .A2(m[8]), .ZN(n_5_2637));
   OAI211_X1 i_5_2986 (.A(n_5_2639), .B(n_5_2642), .C1(n_49), .C2(m[11]), 
      .ZN(n_5_2638));
   NOR2_X1 i_5_2987 (.A1(n_5_2652), .A2(n_5_2909), .ZN(n_5_2639));
   INV_X1 i_5_2988 (.A(n_64), .ZN(n_5_2640));
   INV_X1 i_5_2989 (.A(m[5]), .ZN(n_5_2641));
   AOI21_X1 i_5_2990 (.A(n_5_2739), .B1(n_5_2716), .B2(n_5_2643), .ZN(n_5_2642));
   INV_X1 i_5_2991 (.A(m[10]), .ZN(n_5_2643));
   INV_X1 i_5_2992 (.A(n_5_2645), .ZN(n_5_2644));
   NAND2_X1 i_5_2993 (.A1(n_50), .A2(m[12]), .ZN(n_5_2645));
   NAND2_X1 i_5_2994 (.A1(n_5_2647), .A2(n_5_2648), .ZN(n_5_2646));
   INV_X1 i_5_2995 (.A(n_50), .ZN(n_5_2647));
   INV_X1 i_5_2996 (.A(m[12]), .ZN(n_5_2648));
   NAND2_X1 i_5_2997 (.A1(n_70), .A2(m[6]), .ZN(n_5_2649));
   OAI21_X1 i_5_2998 (.A(n_5_2703), .B1(n_5_2743), .B2(n_5_2739), .ZN(n_5_2650));
   INV_X1 i_5_2999 (.A(n_5_2704), .ZN(n_5_2651));
   INV_X1 i_5_3000 (.A(n_5_2707), .ZN(n_5_2652));
   NAND3_X1 i_5_3001 (.A1(n_70), .A2(n_5_2659), .A3(m[6]), .ZN(n_5_2653));
   NAND3_X1 i_5_3002 (.A1(n_5_2682), .A2(n_5_2657), .A3(n_5_2655), .ZN(n_5_2654));
   NAND2_X1 i_5_3003 (.A1(n_5_2697), .A2(n_5_2656), .ZN(n_5_2655));
   NAND2_X1 i_5_3004 (.A1(n_64), .A2(m[5]), .ZN(n_5_2656));
   INV_X1 i_5_3005 (.A(n_5_2658), .ZN(n_5_2657));
   NAND2_X1 i_5_3006 (.A1(n_5_2659), .A2(n_5_2784), .ZN(n_5_2658));
   OR2_X1 i_5_3007 (.A1(n_62), .A2(m[7]), .ZN(n_5_2659));
   INV_X1 i_5_3008 (.A(n_5_2706), .ZN(n_5_2660));
   INV_X1 i_5_3009 (.A(n_5_2912), .ZN(n_5_2661));
   NOR2_X1 i_5_3010 (.A1(n_77), .A2(m[10]), .ZN(n_5_2662));
   BUF_X1 rt_shieldBuf__2__2__8 (.A(n_5_2629), .Z(n_5_2663));
   NAND2_X1 i_5_3011 (.A1(n_5_2653), .A2(n_5_2609), .ZN(n_5_2664));
   INV_X1 i_5_3012 (.A(n_5_2664), .ZN(n_5_2665));
   NAND2_X1 i_5_3013 (.A1(n_5_2660), .A2(n_5_2703), .ZN(n_5_2666));
   INV_X1 i_5_3014 (.A(n_5_2666), .ZN(n_5_2667));
   NAND2_X1 i_5_3015 (.A1(m[0]), .A2(m[1]), .ZN(n_5_2668));
   INV_X1 i_5_3016 (.A(n_5_2668), .ZN(n_5_2669));
   NAND2_X1 i_5_3017 (.A1(n_5_2735), .A2(n_5_2732), .ZN(n_5_2670));
   INV_X1 i_5_3018 (.A(n_5_2670), .ZN(n_5_2671));
   NAND2_X1 i_5_3019 (.A1(n_72), .A2(m[2]), .ZN(n_5_2672));
   INV_X1 i_5_3020 (.A(n_5_2672), .ZN(n_5_2673));
   NAND2_X1 i_5_3021 (.A1(n_71), .A2(m[3]), .ZN(n_5_2674));
   NOR2_X1 i_5_3022 (.A1(n_5_2669), .A2(m[0]), .ZN(n_5_2675));
   INV_X1 i_5_3023 (.A(n_5_2675), .ZN(n_5_2676));
   NAND3_X1 i_5_3024 (.A1(n_57), .A2(n_63), .A3(n_5_2676), .ZN(n_5_2677));
   INV_X1 i_5_3025 (.A(n_5_2669), .ZN(n_5_2678));
   NOR2_X1 i_5_3026 (.A1(n_5_2675), .A2(n_5_2678), .ZN(n_5_2679));
   NAND2_X1 i_5_3027 (.A1(n_57), .A2(n_5_2679), .ZN(n_5_2680));
   NAND2_X1 i_5_3028 (.A1(n_63), .A2(m[1]), .ZN(n_5_2681));
   OR2_X1 i_5_3029 (.A1(n_70), .A2(m[6]), .ZN(n_5_2682));
   NOR2_X1 i_5_3030 (.A1(n_70), .A2(m[6]), .ZN(n_5_2683));
   AOI21_X1 i_5_3031 (.A(n_5_2683), .B1(n_5_2649), .B2(n_5_2608), .ZN(n_5_2684));
   AOI21_X1 i_5_3032 (.A(n_5_2608), .B1(n_5_2750), .B2(n_5_2656), .ZN(n_5_2685));
   INV_X1 i_5_3033 (.A(n_5_2607), .ZN(n_5_2686));
   NAND2_X1 i_5_3034 (.A1(n_5_2764), .A2(n_5_2686), .ZN(n_5_2687));
   XNOR2_X1 i_5_3035 (.A(n_5_2684), .B(n_5_2686), .ZN(n_5_2688));
   OAI21_X1 i_5_3036 (.A(n_5_2687), .B1(n_5_2688), .B2(n_5_2764), .ZN(n_5_2689));
   NOR2_X1 i_5_3037 (.A1(n_51), .A2(m[13]), .ZN(n_5_2690));
   INV_X1 i_5_3038 (.A(n_51), .ZN(n_5_2691));
   INV_X1 i_5_3039 (.A(m[13]), .ZN(n_5_2692));
   NAND2_X1 i_5_3040 (.A1(n_5_2691), .A2(n_5_2692), .ZN(n_5_2693));
   XNOR2_X1 i_5_3041 (.A(n_67), .B(m[4]), .ZN(n_5_2694));
   NAND3_X1 i_5_3042 (.A1(n_5_2677), .A2(n_5_2680), .A3(n_5_2681), .ZN(n_5_2695));
   NAND3_X1 i_5_3043 (.A1(n_5_2677), .A2(n_5_2680), .A3(n_5_2681), .ZN(n_5_2696));
   NAND2_X1 i_5_3044 (.A1(n_67), .A2(m[4]), .ZN(n_5_2697));
   NAND2_X1 i_5_3045 (.A1(n_67), .A2(m[4]), .ZN(n_5_2698));
   NAND2_X1 i_5_3046 (.A1(n_5_2701), .A2(n_5_2749), .ZN(n_5_2700));
   NAND2_X1 i_5_3047 (.A1(n_5_2650), .A2(n_5_2702), .ZN(n_5_2701));
   NAND2_X1 i_5_3048 (.A1(n_5_2705), .A2(n_5_2704), .ZN(n_5_2702));
   NAND2_X1 i_5_3049 (.A1(n_74), .A2(m[9]), .ZN(n_5_2703));
   NAND2_X1 i_5_3050 (.A1(n_77), .A2(m[10]), .ZN(n_5_2704));
   NAND2_X1 i_5_3051 (.A1(n_5_2716), .A2(n_5_2643), .ZN(n_5_2705));
   INV_X1 i_5_3052 (.A(n_5_2637), .ZN(n_5_2706));
   NAND3_X1 i_5_3053 (.A1(n_5_2776), .A2(n_5_2654), .A3(n_5_2665), .ZN(n_5_2707));
   NAND4_X1 i_5_3054 (.A1(n_5_2776), .A2(n_5_2665), .A3(n_5_2654), .A4(n_5_2637), 
      .ZN(n_5_2708));
   NAND2_X1 i_5_3055 (.A1(n_5_2637), .A2(n_5_2909), .ZN(n_5_2709));
   INV_X1 i_5_3056 (.A(n_5_2723), .ZN(n_5_2710));
   NOR2_X1 i_5_3057 (.A1(n_49), .A2(m[11]), .ZN(n_5_2711));
   INV_X1 i_5_3058 (.A(n_49), .ZN(n_5_2712));
   INV_X1 i_5_3059 (.A(m[11]), .ZN(n_5_2713));
   NAND2_X1 i_5_3060 (.A1(n_5_2712), .A2(n_5_2713), .ZN(n_5_2714));
   AOI21_X1 i_5_3061 (.A(n_5_2745), .B1(n_5_2769), .B2(n_5_2674), .ZN(n_5_2715));
   INV_X1 i_5_3062 (.A(n_77), .ZN(n_5_2716));
   INV_X1 i_5_3063 (.A(n_77), .ZN(n_5_2717));
   INV_X1 i_5_3064 (.A(m[10]), .ZN(n_5_2718));
   INV_X1 i_5_3065 (.A(n_5_2643), .ZN(n_5_2719));
   OAI22_X1 i_5_3066 (.A1(n_5_2717), .A2(n_5_2718), .B1(n_77), .B2(n_5_2719), 
      .ZN(n_5_2720));
   OR2_X1 i_5_3067 (.A1(n_72), .A2(m[2]), .ZN(n_5_2721));
   XNOR2_X1 i_5_3068 (.A(n_72), .B(m[2]), .ZN(n_5_2722));
   NAND2_X1 i_5_3069 (.A1(n_49), .A2(m[11]), .ZN(n_5_2723));
   NAND2_X1 i_5_3070 (.A1(n_5_2662), .A2(m[11]), .ZN(n_5_2724));
   INV_X1 i_5_3071 (.A(n_5_2724), .ZN(n_5_2725));
   NAND2_X1 i_5_3072 (.A1(n_49), .A2(n_5_2725), .ZN(n_5_2726));
   INV_X1 i_5_3073 (.A(n_5_2662), .ZN(n_5_2727));
   OAI21_X1 i_5_3074 (.A(n_5_2726), .B1(n_5_2714), .B2(n_5_2727), .ZN(n_5_2728));
   INV_X1 i_5_3075 (.A(n_5_2704), .ZN(n_5_2729));
   NAND2_X1 i_5_3076 (.A1(n_49), .A2(m[11]), .ZN(n_5_2730));
   AOI21_X1 i_5_3077 (.A(n_5_2729), .B1(n_5_2714), .B2(n_5_2730), .ZN(n_5_2731));
   AOI21_X1 i_5_3078 (.A(n_5_2728), .B1(n_5_2862), .B2(n_5_2731), .ZN(n_5_2732));
   NAND2_X1 i_5_3079 (.A1(n_5_2862), .A2(n_5_2704), .ZN(n_5_2733));
   NOR3_X1 i_5_3080 (.A1(n_5_2710), .A2(n_5_2711), .A3(n_5_2662), .ZN(n_5_2734));
   NAND2_X1 i_5_3081 (.A1(n_5_2733), .A2(n_5_2734), .ZN(n_5_2735));
   NOR2_X1 i_5_3082 (.A1(n_5_2715), .A2(n_5_2752), .ZN(n_5_2736));
   NAND3_X1 i_5_3083 (.A1(n_5_2736), .A2(n_5_2784), .A3(n_5_2656), .ZN(n_5_2737));
   OAI21_X1 i_5_3084 (.A(n_5_2737), .B1(n_5_2788), .B2(n_5_2736), .ZN(n_5_2738));
   NOR2_X1 i_5_3085 (.A1(n_74), .A2(m[9]), .ZN(n_5_2739));
   INV_X1 i_5_3086 (.A(n_74), .ZN(n_5_2740));
   INV_X1 i_5_3087 (.A(m[9]), .ZN(n_5_2741));
   NAND2_X1 i_5_3088 (.A1(n_5_2740), .A2(n_5_2741), .ZN(n_5_2742));
   NAND2_X1 i_5_3089 (.A1(n_5_2708), .A2(n_5_2709), .ZN(n_5_2743));
   NAND2_X1 i_5_3090 (.A1(n_5_2708), .A2(n_5_2709), .ZN(n_5_2744));
   NOR2_X1 i_5_3091 (.A1(n_71), .A2(m[3]), .ZN(n_5_2745));
   INV_X1 i_5_3092 (.A(n_5_2720), .ZN(n_5_2746));
   NAND2_X1 i_5_3093 (.A1(n_5_2703), .A2(n_5_2746), .ZN(n_5_2747));
   INV_X1 i_5_3094 (.A(n_5_2747), .ZN(n_5_2748));
   OAI21_X1 i_5_3095 (.A(n_5_2748), .B1(n_5_2744), .B2(n_5_2739), .ZN(n_5_2749));
   OAI21_X1 i_5_3096 (.A(n_5_2751), .B1(n_5_2771), .B2(n_5_2752), .ZN(n_5_2750));
   OR2_X1 i_5_3097 (.A1(n_67), .A2(m[4]), .ZN(n_5_2751));
   INV_X1 i_5_3098 (.A(n_5_2698), .ZN(n_5_2752));
   NAND2_X1 i_5_3099 (.A1(n_5_2656), .A2(n_5_2674), .ZN(n_5_2753));
   INV_X1 i_5_3100 (.A(n_5_2753), .ZN(n_5_2754));
   INV_X1 i_5_3101 (.A(n_5_2770), .ZN(n_5_2755));
   NAND2_X1 i_5_3102 (.A1(n_5_2755), .A2(n_5_2649), .ZN(n_5_2756));
   NOR2_X1 i_5_3103 (.A1(n_67), .A2(m[4]), .ZN(n_5_2757));
   NAND2_X1 i_5_3104 (.A1(n_5_2656), .A2(n_5_2757), .ZN(n_5_2758));
   INV_X1 i_5_3105 (.A(n_5_2758), .ZN(n_5_2759));
   NAND2_X1 i_5_3106 (.A1(n_5_2649), .A2(n_5_2759), .ZN(n_5_2760));
   NAND3_X1 i_5_3107 (.A1(n_5_2698), .A2(n_5_2656), .A3(n_5_2745), .ZN(n_5_2761));
   INV_X1 i_5_3108 (.A(n_5_2761), .ZN(n_5_2762));
   NAND2_X1 i_5_3109 (.A1(n_5_2649), .A2(n_5_2762), .ZN(n_5_2763));
   NAND3_X1 i_5_3110 (.A1(n_5_2756), .A2(n_5_2760), .A3(n_5_2763), .ZN(n_5_2764));
   NAND3_X1 i_5_3111 (.A1(n_5_2776), .A2(n_5_2665), .A3(n_5_2654), .ZN(n_5_2765));
   NAND2_X1 i_5_3112 (.A1(n_5_2912), .A2(n_5_2637), .ZN(n_5_2766));
   XNOR2_X1 i_5_3113 (.A(n_5_2765), .B(n_5_2766), .ZN(n_5_2767));
   OAI21_X1 i_5_3114 (.A(n_5_2721), .B1(n_5_2696), .B2(n_5_2673), .ZN(n_5_2768));
   OAI21_X1 i_5_3115 (.A(n_5_2721), .B1(n_5_2696), .B2(n_5_2673), .ZN(n_5_2769));
   NAND3_X1 i_5_3116 (.A1(n_5_2769), .A2(n_5_2698), .A3(n_5_2754), .ZN(n_5_2770));
   AOI21_X1 i_5_3117 (.A(n_5_2745), .B1(n_5_2768), .B2(n_5_2674), .ZN(n_5_2771));
   INV_X1 i_5_3118 (.A(m[3]), .ZN(n_5_2772));
   NOR2_X1 i_5_3119 (.A1(n_5_2695), .A2(n_5_2673), .ZN(n_5_2773));
   NAND2_X1 i_5_3120 (.A1(n_5_2783), .A2(n_5_2773), .ZN(n_5_2774));
   OAI21_X1 i_5_3121 (.A(n_5_2774), .B1(n_5_2782), .B2(n_5_2773), .ZN(n_5_2775));
   NAND4_X1 i_5_3122 (.A1(n_5_2682), .A2(n_5_2657), .A3(n_5_2751), .A4(n_5_2778), 
      .ZN(n_5_2776));
   OAI21_X1 i_5_3123 (.A(n_5_2721), .B1(n_5_2695), .B2(n_5_2673), .ZN(n_5_2777));
   AOI21_X1 i_5_3124 (.A(n_5_2745), .B1(n_5_2780), .B2(n_5_2674), .ZN(n_5_2778));
   AOI21_X1 i_5_3125 (.A(n_5_2745), .B1(n_5_2777), .B2(n_5_2674), .ZN(n_5_2779));
   OAI21_X1 i_5_3126 (.A(n_5_2721), .B1(n_5_2695), .B2(n_5_2673), .ZN(n_5_2780));
   XNOR2_X1 i_5_3127 (.A(n_71), .B(n_5_2772), .ZN(n_5_2781));
   XNOR2_X1 i_5_3128 (.A(n_5_2781), .B(n_5_2721), .ZN(n_5_2782));
   XNOR2_X1 i_5_3129 (.A(n_71), .B(n_5_2772), .ZN(n_5_2783));
   NAND2_X1 i_5_3130 (.A1(n_5_2640), .A2(n_5_2641), .ZN(n_5_2784));
   NAND2_X1 i_5_3131 (.A1(n_5_2640), .A2(n_5_2641), .ZN(n_5_2785));
   NAND2_X1 i_5_3132 (.A1(n_5_2656), .A2(n_5_2785), .ZN(n_5_2786));
   INV_X1 i_5_3133 (.A(n_5_2751), .ZN(n_5_2787));
   XNOR2_X1 i_5_3134 (.A(n_5_2786), .B(n_5_2787), .ZN(n_5_2788));
   NAND2_X1 i_5_3135 (.A1(n_5_3008), .A2(m[3]), .ZN(n_5_2789));
   XNOR2_X1 i_5_3136 (.A(n_5_3008), .B(n_5_1892), .ZN(n_5_2790));
   NOR2_X1 i_5_3137 (.A1(n_5_3008), .A2(m[3]), .ZN(n_5_2791));
   XNOR2_X1 i_5_3138 (.A(n_5_3008), .B(n_5_2569), .ZN(n_5_2792));
   NAND2_X1 i_5_3139 (.A1(n_5_3008), .A2(n_5_2569), .ZN(n_5_2793));
   OR2_X1 i_5_3140 (.A1(n_5_3008), .A2(n_5_2569), .ZN(n_5_2794));
   NAND3_X1 i_5_3141 (.A1(n_5_2890), .A2(n_5_2891), .A3(n_5_2358), .ZN(n_5_2795));
   NAND3_X1 i_5_3142 (.A1(n_5_2320), .A2(n_5_2321), .A3(n_5_2322), .ZN(n_5_2796));
   NOR2_X1 i_5_3143 (.A1(n_5_2796), .A2(m[5]), .ZN(n_5_2797));
   XNOR2_X1 i_5_3144 (.A(n_5_2796), .B(n_5_1965), .ZN(n_5_2798));
   NAND2_X1 i_5_3145 (.A1(n_5_2796), .A2(m[5]), .ZN(n_5_2799));
   NAND2_X1 i_5_3146 (.A1(n_5_2803), .A2(n_5_1926), .ZN(n_5_2800));
   XNOR2_X1 i_5_3147 (.A(n_5_2803), .B(n_5_2020), .ZN(n_5_2801));
   NOR2_X1 i_5_3148 (.A1(n_5_2796), .A2(n_66), .ZN(n_5_2802));
   NAND3_X1 i_5_3149 (.A1(n_5_2320), .A2(n_5_2321), .A3(n_5_2322), .ZN(n_5_2803));
   NAND3_X1 i_5_3150 (.A1(n_5_2868), .A2(n_5_2869), .A3(n_5_2360), .ZN(n_5_2804));
   NAND2_X1 i_5_3151 (.A1(n_5_2804), .A2(m[2]), .ZN(n_5_2805));
   NOR2_X1 i_5_3152 (.A1(n_5_2804), .A2(n_5_3329), .ZN(n_5_2806));
   INV_X1 i_5_3153 (.A(n_5_3130), .ZN(n_5_2807));
   NAND3_X1 i_5_3154 (.A1(n_5_2575), .A2(n_5_2576), .A3(n_5_2319), .ZN(n_5_2808));
   XNOR2_X1 i_5_3155 (.A(n_5_2808), .B(n_5_2579), .ZN(n_5_2809));
   NAND2_X1 i_5_3156 (.A1(n_5_2808), .A2(m[4]), .ZN(n_5_2810));
   NAND2_X1 i_5_3157 (.A1(n_5_2808), .A2(m[4]), .ZN(n_5_2811));
   NAND3_X1 i_5_3158 (.A1(n_5_2575), .A2(n_5_2576), .A3(n_5_2319), .ZN(n_5_2812));
   INV_X1 i_5_3159 (.A(n_5_1848), .ZN(n_5_2813));
   INV_X1 i_5_3160 (.A(n_5_1839), .ZN(n_5_2814));
   OAI21_X1 i_5_3161 (.A(n_5_2036), .B1(n_5_2813), .B2(n_5_2814), .ZN(n_5_2815));
   NAND2_X1 i_5_3162 (.A1(n_5_2841), .A2(n_5_2587), .ZN(n_5_2816));
   INV_X1 i_5_3163 (.A(n_5_2816), .ZN(n_5_2817));
   NAND2_X1 i_5_3164 (.A1(n_5_2406), .A2(n_5_2496), .ZN(n_5_2818));
   INV_X1 i_5_3165 (.A(n_5_2818), .ZN(n_5_4078));
   NAND2_X1 i_5_3166 (.A1(n_5_2848), .A2(n_5_4220), .ZN(n_5_2819));
   NAND2_X1 i_5_3167 (.A1(n_5_2323), .A2(n_5_2326), .ZN(n_5_2820));
   NAND2_X1 i_5_3168 (.A1(n_5_2820), .A2(n_5_3185), .ZN(n_5_2821));
   OR2_X1 i_5_3169 (.A1(n_5_2820), .A2(n_5_3185), .ZN(n_5_2822));
   XNOR2_X1 i_5_3170 (.A(n_5_2820), .B(n_5_2145), .ZN(n_5_2823));
   NAND2_X1 i_5_3171 (.A1(n_5_2323), .A2(n_5_2326), .ZN(n_5_2824));
   NAND2_X1 i_5_3172 (.A1(n_5_2602), .A2(n_5_2352), .ZN(n_5_2825));
   INV_X1 i_5_3173 (.A(n_5_2842), .ZN(n_5_2826));
   NAND2_X1 i_5_3174 (.A1(n_5_2524), .A2(n_5_2525), .ZN(n_5_2827));
   INV_X1 i_5_3175 (.A(n_5_2416), .ZN(n_5_2828));
   NAND2_X1 i_5_3176 (.A1(n_5_1927), .A2(n_5_1914), .ZN(n_5_2829));
   INV_X1 i_5_3177 (.A(n_5_2829), .ZN(n_5_2830));
   NOR2_X1 i_5_3178 (.A1(n_5_2824), .A2(m[6]), .ZN(n_5_2831));
   OAI21_X1 i_5_3179 (.A(n_5_2570), .B1(n_5_2824), .B2(m[6]), .ZN(n_5_2832));
   NAND2_X1 i_5_3180 (.A1(n_5_2824), .A2(m[7]), .ZN(n_5_2833));
   NAND2_X1 i_5_3181 (.A1(m[7]), .A2(m[6]), .ZN(n_5_2834));
   XNOR2_X1 i_5_3182 (.A(r[1]), .B(r[0]), .ZN(n_5_2835));
   XNOR2_X1 i_5_3183 (.A(r[1]), .B(r[0]), .ZN(n_5_2836));
   NAND2_X1 i_5_3184 (.A1(n_5_2836), .A2(n_63), .ZN(n_5_2837));
   NAND2_X1 i_5_3185 (.A1(n_5_2356), .A2(n_72), .ZN(n_5_2838));
   INV_X1 i_5_3186 (.A(n_74), .ZN(n_5_2839));
   INV_X1 i_5_3187 (.A(n_74), .ZN(n_5_2840));
   NAND2_X1 i_5_3188 (.A1(n_5_2840), .A2(n_5_2383), .ZN(n_5_2841));
   NAND2_X1 i_5_3189 (.A1(n_5_2542), .A2(n_5_2460), .ZN(n_5_2842));
   NAND2_X1 i_5_3190 (.A1(n_5_2460), .A2(n_5_2542), .ZN(n_5_2843));
   OAI21_X1 i_5_3191 (.A(n_5_2453), .B1(n_5_2454), .B2(n_72), .ZN(n_5_2844));
   INV_X1 i_5_3192 (.A(n_5_2844), .ZN(n_5_4079));
   INV_X1 i_5_3193 (.A(n_5_2405), .ZN(n_5_2845));
   INV_X1 i_5_3194 (.A(n_5_2373), .ZN(n_5_2846));
   AOI21_X1 i_5_3195 (.A(n_5_2846), .B1(n_49), .B2(n_76), .ZN(n_5_2847));
   NAND2_X1 i_5_3196 (.A1(n_5_2845), .A2(n_5_2847), .ZN(n_5_2848));
   NAND2_X1 i_5_3197 (.A1(n_5_2703), .A2(n_5_2742), .ZN(n_5_2849));
   INV_X1 i_5_3198 (.A(n_5_2849), .ZN(n_5_2850));
   NAND2_X1 i_5_3199 (.A1(n_5_2587), .A2(n_5_2359), .ZN(n_5_2851));
   INV_X1 i_5_3200 (.A(n_5_2851), .ZN(n_5_2852));
   NAND2_X1 i_5_3201 (.A1(n_5_2400), .A2(n_5_2852), .ZN(n_5_2853));
   INV_X1 i_5_3202 (.A(n_5_2853), .ZN(n_5_2854));
   NAND2_X1 i_5_3203 (.A1(n_5_2403), .A2(n_5_2359), .ZN(n_5_2855));
   INV_X1 i_5_3204 (.A(n_5_2855), .ZN(n_5_2856));
   INV_X1 i_5_3205 (.A(n_5_2667), .ZN(n_5_2857));
   NOR2_X1 i_5_3206 (.A1(n_74), .A2(m[9]), .ZN(n_5_2858));
   INV_X1 i_5_3207 (.A(n_5_2858), .ZN(n_5_2859));
   INV_X1 i_5_3208 (.A(n_5_2652), .ZN(n_5_2860));
   NOR2_X1 i_5_3209 (.A1(n_5_2661), .A2(n_5_2858), .ZN(n_5_2861));
   AOI22_X1 i_5_3210 (.A1(n_5_2857), .A2(n_5_2859), .B1(n_5_2860), .B2(n_5_2861), 
      .ZN(n_5_2862));
   NAND2_X1 i_5_3211 (.A1(n_5_2352), .A2(n_5_2599), .ZN(n_5_2863));
   NAND2_X1 i_5_3212 (.A1(n_5_4209), .A2(n_5_2361), .ZN(n_5_2864));
   NAND3_X1 i_5_3213 (.A1(n_5_2863), .A2(n_5_2864), .A3(n_5_2837), .ZN(n_5_2865));
   BUF_X1 rt_shieldBuf__2__2__9 (.A(n_69), .Z(n_5_2866));
   NAND3_X1 i_5_3214 (.A1(n_5_2868), .A2(n_5_2869), .A3(n_5_2360), .ZN(n_5_2867));
   NAND2_X1 i_5_3215 (.A1(n_5_2479), .A2(n_5_4209), .ZN(n_5_2868));
   NAND2_X1 i_5_3216 (.A1(n_5_2775), .A2(n_5_2352), .ZN(n_5_2869));
   NAND2_X1 i_5_3217 (.A1(n_5_2479), .A2(n_5_4209), .ZN(n_5_2870));
   NAND2_X1 i_5_3218 (.A1(n_5_2775), .A2(n_5_2352), .ZN(n_5_2871));
   NAND3_X1 i_5_3219 (.A1(n_5_2870), .A2(n_5_2871), .A3(n_5_2360), .ZN(n_5_2872));
   INV_X1 i_5_3220 (.A(n_5_2872), .ZN(n_5_2873));
   NAND3_X1 i_5_3221 (.A1(n_5_2521), .A2(n_5_2592), .A3(n_5_4209), .ZN(n_5_2874));
   NAND2_X1 i_5_3222 (.A1(n_5_2468), .A2(n_5_2520), .ZN(n_5_2875));
   NAND2_X1 i_5_3223 (.A1(n_5_3155), .A2(n_5_2875), .ZN(n_5_2876));
   NAND2_X1 i_5_3224 (.A1(n_5_2889), .A2(n_5_1921), .ZN(n_5_2877));
   NAND2_X1 i_5_3225 (.A1(n_5_1975), .A2(n_5_2080), .ZN(n_5_2878));
   NAND3_X1 i_5_3226 (.A1(n_5_2832), .A2(n_5_2833), .A3(n_5_2834), .ZN(n_5_2879));
   NAND2_X1 i_5_3227 (.A1(n_5_1975), .A2(n_5_2080), .ZN(n_5_2880));
   NAND2_X1 i_5_3228 (.A1(n_5_2889), .A2(n_5_1921), .ZN(n_5_2881));
   NAND3_X1 i_5_3229 (.A1(n_5_2832), .A2(n_5_2833), .A3(n_5_2834), .ZN(n_5_2882));
   NAND3_X1 i_5_3230 (.A1(n_5_2880), .A2(n_5_2881), .A3(n_5_2882), .ZN(n_5_2883));
   XNOR2_X1 i_5_3231 (.A(n_5_2696), .B(n_5_2722), .ZN(n_5_2884));
   NAND2_X1 i_5_3232 (.A1(n_5_2884), .A2(n_5_2352), .ZN(n_5_2885));
   NAND3_X1 i_5_3233 (.A1(n_5_4212), .A2(n_5_2885), .A3(n_5_2838), .ZN(n_5_2886));
   NAND3_X1 i_5_3234 (.A1(n_5_1934), .A2(n_5_1912), .A3(n_5_1913), .ZN(n_5_2887));
   INV_X1 i_5_3235 (.A(n_5_2797), .ZN(n_5_2888));
   NAND2_X1 i_5_3236 (.A1(n_5_2887), .A2(n_5_2888), .ZN(n_5_2889));
   NAND2_X1 i_5_3237 (.A1(n_5_2892), .A2(n_5_4209), .ZN(n_5_2890));
   NAND2_X1 i_5_3238 (.A1(n_5_2893), .A2(n_5_2352), .ZN(n_5_2891));
   XNOR2_X1 i_5_3239 (.A(n_5_2908), .B(n_5_2458), .ZN(n_5_2892));
   XNOR2_X1 i_5_3240 (.A(n_5_2779), .B(n_5_2694), .ZN(n_5_2893));
   XNOR2_X1 i_5_3241 (.A(n_5_2908), .B(n_5_2458), .ZN(n_5_2894));
   XNOR2_X1 i_5_3242 (.A(n_5_2779), .B(n_5_2694), .ZN(n_5_2895));
   NAND3_X1 i_5_3243 (.A1(n_5_2874), .A2(n_5_2825), .A3(n_5_2330), .ZN(n_5_2896));
   NAND2_X1 i_5_3244 (.A1(n_5_2874), .A2(n_5_2330), .ZN(n_5_2897));
   INV_X1 i_5_3245 (.A(n_5_2897), .ZN(n_5_2898));
   NAND2_X1 i_5_3246 (.A1(n_5_2825), .A2(n_5_2898), .ZN(n_5_2899));
   INV_X1 i_5_1682 (.A(n_5_2899), .ZN(n_5_2900));
   NOR2_X1 i_5_3248 (.A1(n_71), .A2(n_65), .ZN(n_5_2901));
   NAND2_X1 i_5_3249 (.A1(n_5_2507), .A2(n_5_2549), .ZN(n_5_2902));
   INV_X1 i_5_3250 (.A(n_71), .ZN(n_5_2903));
   INV_X1 i_5_3251 (.A(n_65), .ZN(n_5_2904));
   NAND2_X1 i_5_3252 (.A1(n_5_2903), .A2(n_5_2904), .ZN(n_5_2905));
   NAND3_X1 i_5_3253 (.A1(n_5_2507), .A2(n_5_2549), .A3(n_5_2905), .ZN(n_5_2906));
   NAND2_X1 i_5_3254 (.A1(n_5_2469), .A2(n_5_2905), .ZN(n_5_2907));
   NAND2_X1 i_5_3255 (.A1(n_5_2906), .A2(n_5_2907), .ZN(n_5_2908));
   NOR2_X1 i_5_3256 (.A1(n_48), .A2(m[8]), .ZN(n_5_2909));
   INV_X1 i_5_3257 (.A(n_48), .ZN(n_5_2910));
   INV_X1 i_5_3258 (.A(m[8]), .ZN(n_5_2911));
   NAND2_X1 i_5_3259 (.A1(n_5_2910), .A2(n_5_2911), .ZN(n_5_2912));
   NAND3_X1 i_5_3260 (.A1(n_5_1829), .A2(n_5_1830), .A3(n_5_1813), .ZN(n_5_2913));
   XNOR2_X1 i_5_3261 (.A(n_5_2913), .B(n_5_2569), .ZN(n_5_2914));
   NAND2_X1 i_5_3262 (.A1(n_5_2918), .A2(m[3]), .ZN(n_5_2915));
   OR2_X1 i_5_3263 (.A1(n_5_2913), .A2(m[3]), .ZN(n_5_2916));
   OR2_X1 i_5_3264 (.A1(n_5_2913), .A2(m[3]), .ZN(n_5_2917));
   NAND3_X1 i_5_3265 (.A1(n_5_1829), .A2(n_5_1830), .A3(n_5_1813), .ZN(n_5_2918));
   NAND2_X1 i_5_3266 (.A1(n_5_1804), .A2(n_5_2916), .ZN(n_5_2919));
   NAND2_X1 i_5_3267 (.A1(n_5_3191), .A2(n_61), .ZN(n_5_2920));
   NAND2_X1 i_5_3268 (.A1(n_5_3853), .A2(n_5_1810), .ZN(n_5_2921));
   NAND2_X1 i_5_3269 (.A1(n_5_3191), .A2(n_61), .ZN(n_5_2922));
   INV_X1 i_5_3270 (.A(n_5_1808), .ZN(n_5_2923));
   NAND3_X1 i_5_3271 (.A1(n_5_2921), .A2(n_5_2922), .A3(n_5_2923), .ZN(n_5_2924));
   NAND2_X1 i_5_3272 (.A1(n_5_2920), .A2(n_5_1805), .ZN(n_5_2925));
   INV_X1 i_5_3273 (.A(n_5_2925), .ZN(n_5_4080));
   INV_X1 i_5_3274 (.A(n_53), .ZN(n_5_2926));
   XNOR2_X1 i_5_3275 (.A(n_5_2218), .B(n_5_2926), .ZN(n_5_2927));
   INV_X1 i_5_3276 (.A(n_5_2218), .ZN(n_5_4081));
   INV_X1 i_5_3277 (.A(n_5_3185), .ZN(n_5_2928));
   INV_X1 i_5_3278 (.A(n_5_1803), .ZN(n_5_2929));
   INV_X1 i_5_3279 (.A(m[6]), .ZN(n_5_2930));
   NAND2_X1 i_5_3280 (.A1(n_5_2116), .A2(n_5_2930), .ZN(n_5_2931));
   INV_X1 i_5_3281 (.A(n_5_2931), .ZN(n_5_2932));
   NAND3_X1 i_5_3282 (.A1(n_5_2986), .A2(n_5_1213), .A3(n_5_2932), .ZN(n_5_2933));
   NAND2_X1 i_5_1888 (.A1(n_5_2221), .A2(n_5_1452), .ZN(n_5_2934));
   NAND2_X1 i_5_3284 (.A1(n_5_3292), .A2(n_5_3293), .ZN(n_5_2935));
   INV_X1 i_5_3285 (.A(n_5_2935), .ZN(n_5_2936));
   INV_X1 i_5_3286 (.A(n_5_2025), .ZN(n_5_2937));
   INV_X1 i_5_3287 (.A(n_5_2011), .ZN(n_5_2938));
   NAND3_X1 i_5_3288 (.A1(n_5_3003), .A2(n_5_2004), .A3(n_5_1986), .ZN(n_5_2939));
   NAND2_X1 i_5_3289 (.A1(n_5_2010), .A2(n_5_1967), .ZN(n_5_2940));
   NAND3_X1 i_5_3290 (.A1(n_5_2004), .A2(n_5_3003), .A3(n_5_1986), .ZN(n_5_2941));
   NAND2_X1 i_5_3291 (.A1(n_5_2010), .A2(n_5_1967), .ZN(n_5_2942));
   NAND2_X1 i_5_3292 (.A1(n_5_2941), .A2(n_5_2942), .ZN(n_5_2943));
   NAND2_X1 i_5_3293 (.A1(n_5_2943), .A2(n_5_2011), .ZN(n_5_2944));
   INV_X1 i_5_3294 (.A(n_5_2944), .ZN(n_5_2945));
   NAND2_X1 i_5_3295 (.A1(n_5_2968), .A2(n_5_3170), .ZN(n_5_2946));
   NAND3_X1 i_5_3296 (.A1(n_5_1438), .A2(n_5_1437), .A3(n_5_1439), .ZN(n_5_2947));
   INV_X1 i_5_3297 (.A(n_5_2947), .ZN(n_5_2948));
   NAND2_X1 i_5_3298 (.A1(n_5_3219), .A2(m[13]), .ZN(n_5_2949));
   NAND2_X1 i_5_3299 (.A1(n_5_3219), .A2(m[13]), .ZN(n_5_2950));
   INV_X1 i_5_3300 (.A(n_5_2950), .ZN(n_5_2951));
   INV_X1 i_5_3301 (.A(n_5_1971), .ZN(n_5_2952));
   NAND2_X1 i_5_3302 (.A1(n_5_4069), .A2(n_76), .ZN(n_5_2953));
   INV_X1 i_5_3303 (.A(n_5_2953), .ZN(n_5_2954));
   NAND2_X1 i_5_3304 (.A1(n_5_4070), .A2(n_5_2954), .ZN(n_5_2955));
   INV_X1 i_5_3305 (.A(n_76), .ZN(n_5_2956));
   INV_X1 i_5_3306 (.A(n_5_4068), .ZN(n_5_2957));
   AOI21_X1 i_5_3307 (.A(n_5_2956), .B1(n_5_4067), .B2(n_5_2957), .ZN(n_5_2958));
   INV_X1 i_5_3308 (.A(n_5_4067), .ZN(n_5_2959));
   OAI21_X1 i_5_3309 (.A(n_5_2958), .B1(n_5_4071), .B2(n_5_2959), .ZN(n_5_2960));
   NAND2_X1 i_5_3310 (.A1(n_5_2955), .A2(n_5_2960), .ZN(n_5_2961));
   INV_X1 i_5_3311 (.A(n_5_2961), .ZN(n_5_2962));
   NAND2_X1 i_5_3312 (.A1(n_5_1784), .A2(n_66), .ZN(n_5_2963));
   INV_X1 i_5_3313 (.A(n_5_2022), .ZN(n_5_2964));
   NAND2_X1 i_5_3314 (.A1(n_5_1784), .A2(n_66), .ZN(n_5_2965));
   NAND2_X1 i_5_3315 (.A1(n_5_2964), .A2(n_5_2965), .ZN(n_5_3188));
   INV_X1 i_5_3316 (.A(n_5_1964), .ZN(n_5_2966));
   NAND2_X1 i_5_3317 (.A1(n_5_2966), .A2(n_5_2965), .ZN(n_5_3189));
   INV_X1 i_5_3318 (.A(m[4]), .ZN(n_5_2967));
   XNOR2_X1 i_5_3319 (.A(n_5_3334), .B(n_5_2919), .ZN(n_5_2968));
   NAND2_X1 i_5_3320 (.A1(n_5_3293), .A2(n_5_3292), .ZN(n_5_2969));
   INV_X1 i_5_3321 (.A(n_5_2969), .ZN(n_5_2970));
   NAND3_X1 i_5_3322 (.A1(n_5_3442), .A2(n_5_3488), .A3(n_5_2159), .ZN(n_5_2971));
   NAND2_X1 i_5_3323 (.A1(n_5_2971), .A2(m[11]), .ZN(n_5_2972));
   XNOR2_X1 i_5_3324 (.A(n_5_3168), .B(n_5_1988), .ZN(n_5_2973));
   NAND2_X1 i_5_3325 (.A1(n_5_1969), .A2(n_5_1970), .ZN(n_5_2974));
   XNOR2_X1 i_5_3326 (.A(n_5_3168), .B(n_5_1988), .ZN(n_5_2975));
   INV_X1 i_5_3327 (.A(n_5_1969), .ZN(n_5_2976));
   NAND2_X1 i_5_3328 (.A1(n_5_2975), .A2(n_5_2976), .ZN(n_5_2977));
   INV_X1 i_5_3329 (.A(n_5_1988), .ZN(n_5_2978));
   XNOR2_X1 i_5_3330 (.A(n_5_2978), .B(n_5_1970), .ZN(n_5_2979));
   XNOR2_X1 i_5_3331 (.A(n_5_3168), .B(n_5_2979), .ZN(n_5_2980));
   NAND2_X1 i_5_3332 (.A1(n_5_2980), .A2(n_5_1969), .ZN(n_5_2981));
   NAND2_X1 i_5_1889 (.A1(n_5_2977), .A2(n_5_2981), .ZN(n_5_2982));
   INV_X1 i_5_3334 (.A(n_5_1979), .ZN(n_5_2983));
   XNOR2_X1 i_5_3335 (.A(n_5_1972), .B(n_5_2983), .ZN(n_5_2984));
   XNOR2_X1 i_5_1705 (.A(n_5_1959), .B(n_5_1950), .ZN(n_5_2985));
   NAND2_X1 i_5_1717 (.A1(n_5_2985), .A2(n_5_3386), .ZN(n_5_2986));
   NAND2_X1 i_5_3338 (.A1(n_5_2300), .A2(n_5_2244), .ZN(n_5_2987));
   INV_X1 i_5_3339 (.A(n_5_2987), .ZN(n_5_2988));
   NAND2_X1 i_5_3340 (.A1(n_5_2138), .A2(n_5_2988), .ZN(n_5_2989));
   INV_X1 i_5_3341 (.A(n_5_2989), .ZN(n_5_2990));
   NAND2_X1 i_5_3342 (.A1(n_5_2134), .A2(n_5_2990), .ZN(n_5_2991));
   XNOR2_X1 i_5_3343 (.A(n_5_2000), .B(n_5_2001), .ZN(n_5_2992));
   XNOR2_X1 i_5_1906 (.A(n_5_2001), .B(n_5_2000), .ZN(n_5_2993));
   NAND2_X1 i_5_1920 (.A1(n_5_2993), .A2(n_5_3170), .ZN(n_5_2994));
   NAND2_X1 i_5_2054 (.A1(n_5_1951), .A2(n_5_3386), .ZN(n_5_2995));
   NAND2_X1 i_5_2091 (.A1(n_5_1989), .A2(n_5_3385), .ZN(n_5_2996));
   NAND2_X1 i_5_3348 (.A1(n_5_2998), .A2(n_5_1966), .ZN(n_5_2997));
   INV_X1 i_5_3349 (.A(n_5_2003), .ZN(n_5_2998));
   NAND2_X1 i_5_3350 (.A1(n_5_2006), .A2(m[1]), .ZN(n_5_2999));
   NAND2_X1 i_5_3351 (.A1(n_5_2006), .A2(m[1]), .ZN(n_5_3000));
   INV_X1 i_5_3352 (.A(n_5_3000), .ZN(n_5_3001));
   INV_X1 i_5_3353 (.A(n_5_1966), .ZN(n_5_3002));
   OAI21_X1 i_5_3354 (.A(n_5_3001), .B1(n_5_2003), .B2(n_5_3002), .ZN(n_5_3003));
   INV_X1 i_5_3355 (.A(n_5_2179), .ZN(n_5_3004));
   NOR2_X1 i_5_3356 (.A1(n_5_2233), .A2(n_5_3004), .ZN(n_5_3005));
   NAND2_X1 i_5_3357 (.A1(n_5_2895), .A2(n_5_2352), .ZN(n_5_3006));
   NAND2_X1 i_5_3358 (.A1(n_5_2894), .A2(n_5_4209), .ZN(n_5_3007));
   NAND3_X1 i_5_3359 (.A1(n_5_3006), .A2(n_5_3007), .A3(n_5_2358), .ZN(n_5_3008));
   NAND2_X1 i_5_3360 (.A1(n_5_1751), .A2(m[11]), .ZN(n_5_3009));
   NAND2_X1 i_5_3361 (.A1(n_5_1982), .A2(n_5_1983), .ZN(n_5_3010));
   NOR2_X1 i_5_3362 (.A1(n_5_2014), .A2(n_5_2952), .ZN(n_5_3011));
   INV_X1 i_5_3363 (.A(n_5_2014), .ZN(n_5_3012));
   INV_X1 i_5_3364 (.A(n_5_2952), .ZN(n_5_3013));
   NAND2_X1 i_5_3365 (.A1(n_5_3012), .A2(n_5_3013), .ZN(n_5_3014));
   NAND3_X1 i_5_3366 (.A1(n_5_1983), .A2(n_5_1982), .A3(n_5_3014), .ZN(n_5_3015));
   NAND2_X1 i_5_3367 (.A1(n_5_1751), .A2(m[11]), .ZN(n_5_3016));
   NAND2_X1 i_5_3368 (.A1(n_5_3015), .A2(n_5_3016), .ZN(n_5_3190));
   NAND2_X1 i_5_3369 (.A1(n_5_1258), .A2(n_5_1259), .ZN(n_5_3017));
   NAND2_X1 i_5_3370 (.A1(n_5_1258), .A2(n_5_1259), .ZN(n_5_3018));
   NAND2_X1 i_5_3371 (.A1(n_5_1526), .A2(n_5_3005), .ZN(n_5_3019));
   NAND2_X1 i_5_3372 (.A1(n_5_3361), .A2(n_5_2180), .ZN(n_5_3020));
   NAND2_X1 i_5_3373 (.A1(n_5_3019), .A2(n_5_3020), .ZN(n_5_3021));
   NAND3_X1 i_5_3374 (.A1(n_5_2994), .A2(n_5_2934), .A3(n_5_2191), .ZN(n_5_3022));
   NOR2_X1 i_5_3375 (.A1(n_5_3022), .A2(n_5_1337), .ZN(n_5_3023));
   INV_X1 i_5_3376 (.A(n_5_3022), .ZN(n_5_3024));
   NAND2_X1 i_5_1718 (.A1(n_5_3029), .A2(m[6]), .ZN(n_5_3025));
   NAND2_X1 i_5_3378 (.A1(n_5_3029), .A2(n_5_3185), .ZN(n_5_3026));
   OAI22_X1 i_5_3379 (.A1(n_5_3024), .A2(n_5_2928), .B1(n_5_3029), .B2(n_5_2929), 
      .ZN(n_5_3027));
   NAND2_X1 i_5_2092 (.A1(n_5_3029), .A2(n_5_3185), .ZN(n_5_3028));
   NAND3_X1 i_5_2103 (.A1(n_5_2994), .A2(n_5_2934), .A3(n_5_2191), .ZN(n_5_3029));
   NAND2_X1 i_5_1762 (.A1(n_5_2807), .A2(n_5_2035), .ZN(n_5_3030));
   INV_X1 i_5_3383 (.A(n_5_2067), .ZN(n_5_3031));
   AOI21_X1 i_5_1763 (.A(n_5_3031), .B1(n_5_3130), .B2(n_5_2034), .ZN(n_5_3032));
   NAND2_X1 i_5_1765 (.A1(n_5_3030), .A2(n_5_3032), .ZN(n_5_3033));
   NAND3_X1 i_5_3386 (.A1(n_5_3742), .A2(n_5_3743), .A3(n_5_3384), .ZN(n_5_3034));
   XOR2_X1 i_5_3387 (.A(n_5_3034), .B(n_66), .Z(n_5_3035));
   XNOR2_X1 i_5_3388 (.A(n_5_3034), .B(m[5]), .ZN(n_5_3036));
   NAND3_X1 i_5_2106 (.A1(n_5_3442), .A2(n_5_3488), .A3(n_5_2159), .ZN(n_5_3037));
   NAND2_X1 i_5_2133 (.A1(n_5_3037), .A2(n_76), .ZN(n_5_3038));
   NAND2_X1 i_5_3391 (.A1(n_5_3068), .A2(n_58), .ZN(n_5_3039));
   INV_X1 i_5_3392 (.A(n_5_3039), .ZN(n_5_3040));
   NAND2_X1 i_5_3393 (.A1(n_5_1944), .A2(n_5_3040), .ZN(n_5_3041));
   NAND2_X1 i_5_3394 (.A1(n_5_1960), .A2(n_5_1871), .ZN(n_5_3042));
   NAND3_X1 i_5_3395 (.A1(n_5_3754), .A2(n_5_3042), .A3(n_5_1923), .ZN(n_5_3337));
   OR2_X1 i_5_3396 (.A1(n_5_3068), .A2(m[4]), .ZN(n_5_3043));
   INV_X1 i_5_3397 (.A(m[4]), .ZN(n_5_3044));
   XNOR2_X1 i_5_3398 (.A(n_5_1945), .B(n_5_3287), .ZN(n_5_3045));
   NAND2_X1 i_5_1766 (.A1(n_5_3045), .A2(n_5_1038), .ZN(n_5_3046));
   INV_X1 i_5_3400 (.A(n_5_3385), .ZN(n_5_3047));
   NAND2_X1 i_5_3401 (.A1(n_5_2155), .A2(n_5_3047), .ZN(n_5_3048));
   NOR2_X1 i_5_3402 (.A1(n_5_2185), .A2(n_5_2189), .ZN(n_5_3049));
   NAND2_X1 i_5_3403 (.A1(n_5_2186), .A2(n_5_2155), .ZN(n_5_3050));
   OAI21_X1 i_5_2166 (.A(n_5_3048), .B1(n_5_3049), .B2(n_5_3050), .ZN(n_5_3051));
   INV_X1 i_5_3405 (.A(n_5_3185), .ZN(n_5_3052));
   NAND2_X1 i_5_3406 (.A1(n_5_2116), .A2(n_5_3052), .ZN(n_5_3053));
   INV_X1 i_5_3407 (.A(n_5_3053), .ZN(n_5_3054));
   NAND3_X1 i_5_3408 (.A1(n_5_2049), .A2(n_5_2050), .A3(n_5_2051), .ZN(n_5_3055));
   NOR2_X1 i_5_3409 (.A1(n_5_3055), .A2(n_5_2568), .ZN(n_5_3056));
   NAND2_X1 i_5_3410 (.A1(n_5_3063), .A2(n_5_2568), .ZN(n_5_3057));
   NAND2_X1 i_5_3411 (.A1(n_5_3055), .A2(n_5_2568), .ZN(n_5_3058));
   INV_X1 i_5_3412 (.A(n_5_3063), .ZN(n_5_3059));
   INV_X1 i_5_3413 (.A(n_5_3055), .ZN(n_5_3060));
   NOR2_X1 i_5_3414 (.A1(n_5_3055), .A2(m[1]), .ZN(n_5_3061));
   NAND2_X1 i_5_3415 (.A1(n_5_3055), .A2(m[1]), .ZN(n_5_3062));
   NAND3_X1 i_5_3416 (.A1(n_5_2049), .A2(n_5_2050), .A3(n_5_2051), .ZN(n_5_3063));
   NAND2_X1 i_5_3417 (.A1(n_5_4534), .A2(n_5_1850), .ZN(n_5_3064));
   NAND2_X1 i_5_3418 (.A1(n_5_4534), .A2(n_5_1850), .ZN(n_5_3065));
   NAND2_X1 i_5_3419 (.A1(n_5_678), .A2(m[12]), .ZN(n_5_3066));
   NAND2_X1 i_5_698 (.A1(n_5_3065), .A2(n_5_3066), .ZN(n_5_3067));
   NAND3_X1 i_5_3421 (.A1(n_5_3132), .A2(n_5_3378), .A3(n_5_1212), .ZN(n_5_3068));
   NAND3_X1 i_5_3422 (.A1(n_5_2090), .A2(n_5_3459), .A3(n_5_2110), .ZN(n_5_3069));
   OR2_X1 i_5_3423 (.A1(n_5_3069), .A2(n_65), .ZN(n_5_3397));
   OR2_X1 i_5_3424 (.A1(n_5_3069), .A2(n_65), .ZN(n_5_3070));
   XNOR2_X1 i_5_3425 (.A(n_5_3069), .B(n_65), .ZN(n_5_3071));
   INV_X1 i_5_3426 (.A(n_5_3398), .ZN(n_5_3072));
   OAI21_X1 i_5_3427 (.A(n_5_3072), .B1(n_5_3069), .B2(n_5_2005), .ZN(n_5_3073));
   AOI21_X1 i_5_3428 (.A(n_5_2023), .B1(n_5_3069), .B2(n_5_1999), .ZN(n_5_3074));
   NOR2_X1 i_5_3429 (.A1(n_5_3069), .A2(m[3]), .ZN(n_5_3075));
   NAND2_X1 i_5_3430 (.A1(n_5_3069), .A2(m[3]), .ZN(n_5_3076));
   NAND3_X1 i_5_3431 (.A1(n_5_2090), .A2(n_5_3459), .A3(n_5_2110), .ZN(n_5_3398));
   XNOR2_X1 i_5_1767 (.A(n_5_2267), .B(n_5_3260), .ZN(n_5_3077));
   NAND2_X1 i_5_1812 (.A1(n_5_3077), .A2(n_5_4068), .ZN(n_5_3078));
   NAND2_X1 i_5_3434 (.A1(n_5_1998), .A2(n_5_1036), .ZN(n_5_3079));
   NAND3_X1 i_5_3435 (.A1(n_5_3504), .A2(n_5_3079), .A3(n_5_1938), .ZN(n_5_3399));
   AOI21_X1 i_5_707 (.A(n_5_1826), .B1(n_5_1828), .B2(n_5_1863), .ZN(n_5_3080));
   NAND2_X1 i_5_3437 (.A1(n_5_1828), .A2(n_5_1863), .ZN(n_5_3081));
   INV_X1 i_5_3438 (.A(m[12]), .ZN(n_5_3082));
   NAND2_X1 i_5_3439 (.A1(n_5_4061), .A2(n_5_3082), .ZN(n_5_3083));
   INV_X1 i_5_3440 (.A(n_5_3083), .ZN(n_5_3084));
   NAND3_X1 i_5_3441 (.A1(n_5_4059), .A2(n_5_4060), .A3(n_5_3084), .ZN(n_5_3085));
   INV_X1 i_5_3442 (.A(n_5_3085), .ZN(n_5_3086));
   NOR2_X1 i_5_3443 (.A1(n_5_1826), .A2(n_5_3086), .ZN(n_5_3087));
   NAND2_X1 i_5_3444 (.A1(n_5_3081), .A2(n_5_3087), .ZN(n_5_3088));
   INV_X1 i_5_3445 (.A(n_5_3185), .ZN(n_5_3089));
   NAND2_X1 i_5_3446 (.A1(n_5_2191), .A2(n_5_3089), .ZN(n_5_3090));
   INV_X1 i_5_3447 (.A(n_5_3090), .ZN(n_5_3091));
   NAND3_X1 i_5_3448 (.A1(n_5_3305), .A2(n_5_3306), .A3(n_5_3091), .ZN(n_5_3092));
   INV_X1 i_5_3449 (.A(n_5_3092), .ZN(n_5_3093));
   NAND3_X1 i_5_3450 (.A1(n_5_2251), .A2(n_5_2252), .A3(n_5_2240), .ZN(n_5_3094));
   NAND3_X1 i_5_3451 (.A1(n_5_2251), .A2(n_5_2252), .A3(n_5_2240), .ZN(n_5_3095));
   INV_X1 i_5_3452 (.A(n_5_3095), .ZN(n_5_3096));
   NAND2_X1 i_5_3453 (.A1(n_5_2253), .A2(n_5_4069), .ZN(n_5_3097));
   INV_X1 i_5_3454 (.A(n_5_2248), .ZN(n_5_3098));
   AOI21_X1 i_5_3455 (.A(n_5_3098), .B1(n_5_2262), .B2(n_5_4068), .ZN(n_5_3099));
   NAND2_X1 i_5_3456 (.A1(n_5_3097), .A2(n_5_3099), .ZN(n_5_3191));
   NAND3_X1 i_5_3457 (.A1(n_5_2235), .A2(n_5_2207), .A3(n_5_2210), .ZN(n_5_3100));
   NAND2_X1 i_5_3458 (.A1(n_5_2236), .A2(n_5_2237), .ZN(n_5_3101));
   NAND2_X1 i_5_3459 (.A1(n_5_3100), .A2(n_5_3101), .ZN(n_5_3102));
   NAND2_X1 i_5_3460 (.A1(n_5_2217), .A2(n_5_2214), .ZN(n_5_3103));
   INV_X1 i_5_3461 (.A(n_5_3103), .ZN(n_5_3104));
   NOR2_X1 i_5_2167 (.A1(n_5_2229), .A2(n_5_3093), .ZN(n_5_3105));
   NAND2_X1 i_5_2168 (.A1(n_5_3546), .A2(n_5_3105), .ZN(n_5_3106));
   NAND3_X1 i_5_3464 (.A1(n_5_2241), .A2(n_5_2242), .A3(n_5_2243), .ZN(n_5_3107));
   NAND2_X1 i_5_3465 (.A1(n_5_2242), .A2(n_5_2243), .ZN(n_5_3108));
   INV_X1 i_5_3466 (.A(n_5_3108), .ZN(n_5_3109));
   NAND2_X1 i_5_3467 (.A1(n_5_2241), .A2(n_5_3109), .ZN(n_5_3110));
   INV_X1 i_5_3468 (.A(n_5_3110), .ZN(n_5_3111));
   INV_X1 i_5_2302 (.A(n_5_3093), .ZN(n_5_3112));
   NAND3_X1 i_5_1813 (.A1(n_5_2197), .A2(n_5_2198), .A3(n_5_2192), .ZN(n_5_3113));
   NAND3_X1 i_5_3471 (.A1(n_5_2197), .A2(n_5_2198), .A3(n_5_2192), .ZN(n_5_3114));
   INV_X1 i_5_3472 (.A(n_5_3114), .ZN(n_5_3115));
   INV_X1 i_5_3473 (.A(n_5_3094), .ZN(n_5_3116));
   NAND2_X1 i_5_3474 (.A1(n_5_2208), .A2(n_5_3116), .ZN(n_5_3117));
   INV_X1 i_5_3475 (.A(n_5_2209), .ZN(n_5_3118));
   NAND2_X1 i_5_3476 (.A1(n_5_3117), .A2(n_5_3118), .ZN(n_5_3119));
   INV_X1 i_5_3477 (.A(n_5_2208), .ZN(n_5_3120));
   NAND2_X1 i_5_3478 (.A1(n_5_3120), .A2(n_5_3116), .ZN(n_5_3121));
   NAND2_X1 i_5_3479 (.A1(n_5_3119), .A2(n_5_3121), .ZN(n_5_3122));
   AOI21_X1 i_5_3480 (.A(n_5_2332), .B1(n_5_2438), .B2(n_5_2856), .ZN(n_5_3123));
   NAND2_X1 i_5_3481 (.A1(n_5_2854), .A2(n_5_2445), .ZN(n_5_3125));
   NAND2_X1 i_5_3482 (.A1(n_5_2700), .A2(n_5_2352), .ZN(n_5_3127));
   NAND3_X1 i_5_1846 (.A1(n_5_3123), .A2(n_5_3125), .A3(n_5_3127), .ZN(n_5_3130));
   NAND2_X1 i_5_3484 (.A1(n_5_3236), .A2(n_5_3385), .ZN(n_5_3132));
   AOI21_X1 i_5_3485 (.A(n_5_2212), .B1(n_5_3122), .B2(n_5_2213), .ZN(n_5_3133));
   NAND2_X1 i_5_3333 (.A1(n_5_3234), .A2(n_5_1452), .ZN(n_5_3134));
   AOI21_X1 i_5_3344 (.A(n_5_2212), .B1(n_5_3122), .B2(n_5_2213), .ZN(n_5_3135));
   NAND2_X1 i_5_3345 (.A1(n_5_3134), .A2(n_5_3135), .ZN(n_5_3137));
   NAND3_X1 i_5_3489 (.A1(n_5_3408), .A2(n_5_2088), .A3(n_5_2089), .ZN(n_5_3140));
   INV_X1 i_5_3490 (.A(n_5_3329), .ZN(n_5_3144));
   NAND2_X1 i_5_3491 (.A1(n_5_2089), .A2(n_5_3144), .ZN(n_5_3145));
   INV_X1 i_5_3492 (.A(n_5_3145), .ZN(n_5_3146));
   NAND3_X1 i_5_3493 (.A1(n_5_3408), .A2(n_5_2088), .A3(n_5_3146), .ZN(n_5_3150));
   NAND2_X1 i_5_3494 (.A1(n_5_2524), .A2(n_5_2525), .ZN(n_5_3153));
   NOR2_X1 i_5_3495 (.A1(n_5_2843), .A2(n_5_2416), .ZN(n_5_3154));
   NAND2_X1 i_5_3496 (.A1(n_5_3153), .A2(n_5_3154), .ZN(n_5_3155));
   AND3_X1 i_5_3497 (.A1(n_5_2255), .A2(n_5_2254), .A3(n_5_2256), .ZN(n_5_3156));
   NAND2_X1 i_5_3498 (.A1(n_5_2254), .A2(n_5_2261), .ZN(n_5_3159));
   INV_X1 i_5_3499 (.A(n_5_3159), .ZN(n_5_3161));
   NAND3_X1 i_5_3500 (.A1(n_5_2255), .A2(n_5_2256), .A3(n_5_3161), .ZN(n_5_3169));
   INV_X1 i_5_3501 (.A(n_5_2169), .ZN(n_5_3184));
   NAND2_X1 i_5_3502 (.A1(n_5_3213), .A2(n_5_2219), .ZN(n_5_3186));
   INV_X1 i_5_3503 (.A(n_5_3186), .ZN(n_5_3187));
   XNOR2_X1 i_5_3504 (.A(n_5_2228), .B(m[8]), .ZN(n_5_3192));
   NOR2_X1 i_5_3505 (.A1(n_5_2188), .A2(n_5_2211), .ZN(n_5_3193));
   NAND2_X1 i_5_3506 (.A1(n_5_3192), .A2(n_5_3193), .ZN(n_5_3194));
   XNOR2_X1 i_5_3507 (.A(n_5_2187), .B(m[8]), .ZN(n_5_3195));
   XNOR2_X1 i_5_3508 (.A(n_5_3195), .B(n_5_2228), .ZN(n_5_3196));
   OAI21_X1 i_5_3509 (.A(n_5_3194), .B1(n_5_3196), .B2(n_5_3193), .ZN(n_5_3197));
   NAND2_X1 i_5_3346 (.A1(n_5_3486), .A2(n_5_3385), .ZN(n_5_3198));
   NAND2_X1 i_5_3511 (.A1(n_5_2174), .A2(n_5_3386), .ZN(n_5_4082));
   NAND2_X1 i_5_3512 (.A1(n_5_3197), .A2(n_5_3385), .ZN(n_5_4083));
   NAND2_X1 i_5_3513 (.A1(n_5_3137), .A2(n_5_2165), .ZN(n_5_4084));
   NAND2_X1 i_5_3514 (.A1(n_5_678), .A2(m[12]), .ZN(n_5_3199));
   NAND2_X1 i_5_3515 (.A1(n_5_3080), .A2(n_5_3064), .ZN(n_5_3200));
   NAND2_X1 i_5_3516 (.A1(n_5_678), .A2(m[12]), .ZN(n_5_3201));
   NAND2_X1 i_5_3517 (.A1(n_5_3200), .A2(n_5_3201), .ZN(n_5_3202));
   XNOR2_X1 i_5_3518 (.A(n_5_1734), .B(n_5_1778), .ZN(n_5_3203));
   NAND2_X1 i_5_3381 (.A1(n_5_3203), .A2(n_5_3386), .ZN(n_5_3204));
   NAND2_X1 i_5_3520 (.A1(n_5_1819), .A2(n_5_1806), .ZN(n_5_3205));
   NAND2_X1 i_5_3521 (.A1(n_5_3202), .A2(n_5_1844), .ZN(n_5_3206));
   INV_X1 i_5_3522 (.A(n_5_1820), .ZN(n_5_3207));
   NAND3_X1 i_5_3523 (.A1(n_5_3205), .A2(n_5_3206), .A3(n_5_3207), .ZN(n_5_3208));
   NAND2_X1 i_5_3524 (.A1(n_5_3208), .A2(n_5_1817), .ZN(n_5_3209));
   NAND2_X1 i_5_3525 (.A1(n_5_3180), .A2(n_5_3336), .ZN(n_5_3210));
   INV_X1 i_5_3526 (.A(n_5_3210), .ZN(n_5_3211));
   NAND2_X1 i_5_3527 (.A1(n_5_3181), .A2(n_5_3211), .ZN(n_5_3212));
   INV_X1 i_5_3528 (.A(n_5_3212), .ZN(n_5_3213));
   NAND2_X1 i_5_3529 (.A1(n_5_2202), .A2(n_5_2199), .ZN(n_5_3214));
   NAND3_X1 i_5_3530 (.A1(n_5_3374), .A2(n_5_2204), .A3(n_5_3525), .ZN(n_5_3215));
   NAND2_X1 i_5_3531 (.A1(n_5_3214), .A2(n_5_3215), .ZN(n_5_3216));
   NAND2_X1 i_5_1805 (.A1(n_5_3925), .A2(n_5_3385), .ZN(n_5_3217));
   NAND2_X1 i_5_1806 (.A1(n_5_2168), .A2(n_5_3386), .ZN(n_5_3218));
   NAND3_X1 i_5_2019 (.A1(n_5_3217), .A2(n_5_3218), .A3(n_5_2166), .ZN(n_5_3219));
   NAND2_X1 i_5_3535 (.A1(n_5_2191), .A2(n_5_2181), .ZN(n_5_3220));
   INV_X1 i_5_3536 (.A(n_5_3220), .ZN(n_5_3221));
   NAND3_X1 i_5_3537 (.A1(n_5_3305), .A2(n_5_3306), .A3(n_5_3221), .ZN(n_5_3222));
   NOR2_X1 i_5_3538 (.A1(n_5_2570), .A2(m[7]), .ZN(n_5_3223));
   INV_X1 i_5_3539 (.A(n_5_2570), .ZN(n_5_3224));
   INV_X1 i_5_3540 (.A(m[7]), .ZN(n_5_3225));
   NAND2_X1 i_5_3541 (.A1(n_5_3224), .A2(n_5_3225), .ZN(n_5_3226));
   XNOR2_X1 i_5_3542 (.A(n_5_3457), .B(n_5_2170), .ZN(n_5_3227));
   INV_X1 i_5_3543 (.A(n_5_2866), .ZN(n_5_3228));
   NAND3_X1 i_5_3382 (.A1(n_5_3204), .A2(n_5_3198), .A3(n_5_2159), .ZN(n_5_3229));
   INV_X1 i_5_3545 (.A(m[11]), .ZN(n_5_3230));
   NAND2_X1 i_5_3546 (.A1(n_5_2159), .A2(n_5_3230), .ZN(n_5_3231));
   INV_X1 i_5_3547 (.A(n_5_3231), .ZN(n_5_3232));
   NAND3_X1 i_5_3548 (.A1(n_5_3204), .A2(n_5_3198), .A3(n_5_3232), .ZN(n_5_3233));
   XNOR2_X1 i_5_3549 (.A(n_5_3178), .B(n_5_3179), .ZN(n_5_3234));
   NAND2_X1 i_5_3550 (.A1(n_5_3300), .A2(n_5_1038), .ZN(n_5_3235));
   XNOR2_X1 i_5_3551 (.A(n_5_2182), .B(n_5_2190), .ZN(n_5_3236));
   XNOR2_X1 i_5_3552 (.A(n_5_2182), .B(n_5_2190), .ZN(n_5_3237));
   INV_X1 i_5_3553 (.A(n_5_3239), .ZN(n_5_3238));
   NAND2_X1 i_5_3554 (.A1(n_5_2232), .A2(m[4]), .ZN(n_5_3239));
   NAND2_X1 i_5_3555 (.A1(n_5_2232), .A2(m[4]), .ZN(n_5_3240));
   INV_X1 i_5_3556 (.A(n_5_3240), .ZN(n_5_3241));
   INV_X1 i_5_3557 (.A(n_5_2180), .ZN(n_5_3242));
   OAI21_X1 i_5_3558 (.A(n_5_3241), .B1(n_5_2234), .B2(n_5_3242), .ZN(n_5_3243));
   NAND2_X1 i_5_3559 (.A1(n_5_2270), .A2(n_5_2304), .ZN(n_5_3244));
   INV_X1 i_5_3560 (.A(n_5_3244), .ZN(n_5_3245));
   NAND3_X1 i_5_3561 (.A1(n_5_2245), .A2(n_5_2247), .A3(n_5_2248), .ZN(n_5_3246));
   INV_X1 i_5_3562 (.A(m[14]), .ZN(n_5_3247));
   NAND2_X1 i_5_3563 (.A1(n_5_2248), .A2(n_5_3247), .ZN(n_5_3248));
   INV_X1 i_5_3564 (.A(n_5_3248), .ZN(n_5_3249));
   NAND3_X1 i_5_3565 (.A1(n_5_2245), .A2(n_5_2247), .A3(n_5_3249), .ZN(n_5_4085));
   NAND2_X1 i_5_3566 (.A1(n_5_2811), .A2(n_5_2258), .ZN(n_5_3250));
   INV_X1 i_5_3567 (.A(n_5_3250), .ZN(n_5_3251));
   NAND3_X1 i_5_3568 (.A1(n_5_3251), .A2(n_5_2800), .A3(n_5_2257), .ZN(n_5_3252));
   AOI21_X1 i_5_3569 (.A(n_5_3075), .B1(n_5_2029), .B2(n_5_3076), .ZN(n_5_3253));
   OAI21_X1 i_5_1924 (.A(n_5_3417), .B1(n_5_3472), .B2(n_5_3253), .ZN(n_5_3254));
   NAND2_X1 i_5_3571 (.A1(n_5_3245), .A2(n_5_2269), .ZN(n_5_3255));
   AOI22_X1 i_5_3572 (.A1(n_5_2276), .A2(n_5_2278), .B1(n_5_2304), .B2(n_5_2268), 
      .ZN(n_5_3256));
   INV_X1 i_5_3573 (.A(n_5_2271), .ZN(n_5_3257));
   NAND2_X1 i_5_3574 (.A1(n_5_3245), .A2(n_5_2269), .ZN(n_5_3258));
   AOI22_X1 i_5_3575 (.A1(n_5_2276), .A2(n_5_2278), .B1(n_5_2304), .B2(n_5_2268), 
      .ZN(n_5_3259));
   AOI21_X1 i_5_1950 (.A(n_5_3257), .B1(n_5_3258), .B2(n_5_3259), .ZN(n_5_3260));
   NAND3_X1 i_5_3577 (.A1(n_5_3306), .A2(n_5_3305), .A3(n_5_2191), .ZN(n_5_3261));
   INV_X1 i_5_3578 (.A(n_5_3346), .ZN(n_5_3262));
   NAND2_X1 i_5_3579 (.A1(n_5_3348), .A2(n_58), .ZN(n_5_3263));
   NAND2_X1 i_5_3580 (.A1(n_5_3418), .A2(n_5_3185), .ZN(n_5_3264));
   NAND2_X1 i_5_3581 (.A1(n_5_3746), .A2(n_66), .ZN(n_5_3265));
   NAND2_X1 i_5_3582 (.A1(n_5_2116), .A2(n_5_3384), .ZN(n_5_3266));
   INV_X1 i_5_3583 (.A(n_5_3266), .ZN(n_5_3267));
   NAND3_X1 i_5_3584 (.A1(n_5_3742), .A2(n_5_3743), .A3(n_5_3267), .ZN(n_5_3268));
   INV_X1 i_5_3585 (.A(n_66), .ZN(n_5_3269));
   NAND2_X1 i_5_3586 (.A1(n_5_2116), .A2(n_5_3269), .ZN(n_5_3270));
   INV_X1 i_5_3587 (.A(n_5_3270), .ZN(n_5_3271));
   INV_X1 i_5_3588 (.A(n_5_2116), .ZN(n_5_3272));
   NAND2_X1 i_5_3589 (.A1(n_5_3272), .A2(n_5_3185), .ZN(n_5_3273));
   AOI21_X1 i_5_3590 (.A(n_5_3271), .B1(n_5_3054), .B2(n_5_3273), .ZN(n_5_3274));
   NAND2_X1 i_5_3591 (.A1(n_5_3268), .A2(n_5_3274), .ZN(n_5_3275));
   NAND3_X1 i_5_3592 (.A1(n_5_3275), .A2(n_5_2986), .A3(n_5_1213), .ZN(n_5_3276));
   INV_X1 i_5_3593 (.A(n_5_3185), .ZN(n_5_3277));
   NAND2_X1 i_5_3594 (.A1(n_5_3384), .A2(n_5_3277), .ZN(n_5_3278));
   INV_X1 i_5_3595 (.A(n_5_3278), .ZN(n_5_3279));
   NAND3_X1 i_5_3596 (.A1(n_5_3742), .A2(n_5_3743), .A3(n_5_3279), .ZN(n_5_3280));
   NAND2_X1 i_5_3597 (.A1(n_5_3277), .A2(n_5_3269), .ZN(n_5_3281));
   NAND2_X1 i_5_3598 (.A1(n_5_3280), .A2(n_5_3281), .ZN(n_5_3282));
   INV_X1 i_5_3599 (.A(n_5_3282), .ZN(n_5_3283));
   NAND2_X1 i_5_3600 (.A1(n_5_3276), .A2(n_5_3283), .ZN(n_5_3284));
   NAND3_X1 i_5_3389 (.A1(n_5_2995), .A2(n_5_2996), .A3(n_5_2153), .ZN(n_5_3285));
   NOR2_X1 i_5_3390 (.A1(n_5_3285), .A2(n_60), .ZN(n_5_3286));
   XNOR2_X1 i_5_3603 (.A(n_5_3285), .B(n_60), .ZN(n_5_3287));
   NAND2_X1 i_5_3604 (.A1(n_5_3291), .A2(m[8]), .ZN(n_5_3288));
   OR2_X1 i_5_3605 (.A1(n_5_3285), .A2(m[8]), .ZN(n_5_3289));
   XNOR2_X1 i_5_3606 (.A(n_5_3285), .B(m[8]), .ZN(n_5_3290));
   NAND3_X1 i_5_3420 (.A1(n_5_2995), .A2(n_5_2996), .A3(n_5_2153), .ZN(n_5_3291));
   NAND2_X1 i_5_3608 (.A1(n_5_2216), .A2(n_5_1452), .ZN(n_5_3292));
   AOI21_X1 i_5_3609 (.A(n_5_2196), .B1(n_5_2203), .B2(n_5_3170), .ZN(n_5_3293));
   NAND2_X1 i_5_3610 (.A1(n_5_2203), .A2(n_5_3170), .ZN(n_5_3294));
   NAND2_X1 i_5_3611 (.A1(n_5_2216), .A2(n_5_1452), .ZN(n_5_3295));
   INV_X1 i_5_3612 (.A(n_5_2196), .ZN(n_5_3296));
   NAND3_X1 i_5_3613 (.A1(n_5_3294), .A2(n_5_3295), .A3(n_5_3296), .ZN(n_5_3297));
   INV_X1 i_5_3614 (.A(n_5_1942), .ZN(n_5_3298));
   XNOR2_X1 i_5_3615 (.A(n_5_3140), .B(n_5_3298), .ZN(n_5_3299));
   XNOR2_X1 i_5_3616 (.A(n_5_3299), .B(n_5_1956), .ZN(n_5_3300));
   NAND2_X1 i_5_3617 (.A1(n_5_3435), .A2(n_5_3070), .ZN(n_5_3301));
   NAND2_X1 i_5_3618 (.A1(n_5_3068), .A2(n_58), .ZN(n_5_3302));
   NAND2_X1 i_5_3619 (.A1(n_5_3398), .A2(n_65), .ZN(n_5_3303));
   NAND3_X1 i_5_3620 (.A1(n_5_3301), .A2(n_5_3302), .A3(n_5_3303), .ZN(n_5_3304));
   NAND2_X1 i_5_3621 (.A1(n_5_2992), .A2(n_5_3170), .ZN(n_5_3305));
   NAND2_X1 i_5_3622 (.A1(n_5_2221), .A2(n_5_1452), .ZN(n_5_3306));
   INV_X1 i_5_3623 (.A(n_5_1452), .ZN(n_5_3307));
   NAND2_X1 i_5_3624 (.A1(n_5_2191), .A2(n_5_3307), .ZN(n_5_3308));
   NAND2_X1 i_5_3625 (.A1(n_5_2221), .A2(n_5_3308), .ZN(n_5_3309));
   NAND2_X1 i_5_3626 (.A1(n_5_2992), .A2(n_5_3170), .ZN(n_5_3310));
   INV_X1 i_5_3627 (.A(n_5_2191), .ZN(n_5_3311));
   NAND2_X1 i_5_3628 (.A1(n_5_3308), .A2(n_5_3311), .ZN(n_5_3312));
   NAND3_X1 i_5_3629 (.A1(n_5_3309), .A2(n_5_3310), .A3(n_5_3312), .ZN(n_5_3313));
   INV_X1 i_5_1981 (.A(n_5_3313), .ZN(n_5_3314));
   NAND3_X1 i_5_3631 (.A1(n_5_1074), .A2(n_5_1943), .A3(n_5_3058), .ZN(n_5_3315));
   NAND2_X1 i_5_3632 (.A1(n_5_1968), .A2(n_5_1036), .ZN(n_5_3316));
   NAND3_X1 i_5_1983 (.A1(n_5_3316), .A2(n_5_3791), .A3(n_5_1924), .ZN(n_5_3401));
   NAND3_X1 i_5_3436 (.A1(n_5_2160), .A2(n_5_2161), .A3(n_5_2162), .ZN(n_5_3317));
   INV_X1 i_5_3635 (.A(n_5_3317), .ZN(n_5_3318));
   XNOR2_X1 i_5_3462 (.A(n_5_3317), .B(n_75), .ZN(n_5_3319));
   NAND3_X1 i_5_3463 (.A1(n_5_2160), .A2(n_5_2161), .A3(n_5_2162), .ZN(n_5_3320));
   NAND3_X1 i_5_3638 (.A1(n_5_2265), .A2(n_5_2263), .A3(n_5_2239), .ZN(n_5_3321));
   INV_X1 i_5_3639 (.A(n_5_2264), .ZN(n_5_3322));
   NAND2_X1 i_5_3640 (.A1(n_5_3322), .A2(n_5_4068), .ZN(n_5_3323));
   INV_X1 i_5_3641 (.A(n_5_2239), .ZN(n_5_3324));
   INV_X1 i_5_3642 (.A(n_5_2266), .ZN(n_5_3325));
   AOI21_X1 i_5_3643 (.A(n_5_3324), .B1(n_5_3325), .B2(n_5_4068), .ZN(n_5_3326));
   NAND2_X1 i_5_3644 (.A1(n_5_3323), .A2(n_5_3326), .ZN(n_5_3327));
   NAND2_X1 i_5_3645 (.A1(n_5_3321), .A2(n_5_3327), .ZN(n_5_3328));
   BUF_X1 rt_shieldBuf__2__2__10 (.A(n_59), .Z(n_5_3329));
   NAND4_X1 i_5_3646 (.A1(n_5_3570), .A2(n_5_1953), .A3(n_5_3304), .A4(n_5_1944), 
      .ZN(n_5_3330));
   NAND3_X1 i_5_3647 (.A1(n_5_2249), .A2(n_5_2250), .A3(n_5_2238), .ZN(n_5_3331));
   XNOR2_X1 i_5_3648 (.A(n_5_3348), .B(n_5_2967), .ZN(n_5_3334));
   OR2_X1 i_5_3649 (.A1(n_5_3331), .A2(n_58), .ZN(n_5_3336));
   XNOR2_X1 i_5_3650 (.A(n_5_3331), .B(n_58), .ZN(n_5_3342));
   NAND2_X1 i_5_3651 (.A1(n_5_3331), .A2(m[4]), .ZN(n_5_3344));
   NAND2_X1 i_5_3652 (.A1(n_5_3331), .A2(n_58), .ZN(n_5_3346));
   NAND3_X1 i_5_3653 (.A1(n_5_2249), .A2(n_5_2250), .A3(n_5_2238), .ZN(n_5_3348));
   XNOR2_X1 i_5_3654 (.A(n_5_2259), .B(n_5_2260), .ZN(n_5_3349));
   NAND2_X1 i_5_3655 (.A1(n_5_3349), .A2(n_5_4069), .ZN(n_5_3351));
   MUX2_X1 i_5_3656 (.A(n_5_2218), .B(n_5_2927), .S(n_5_3246), .Z(n_5_3403));
   NAND2_X1 i_5_3469 (.A1(n_5_4174), .A2(n_5_1036), .ZN(n_5_462));
   NAND2_X1 i_5_3658 (.A1(n_5_3361), .A2(n_5_2180), .ZN(n_5_3354));
   NAND2_X1 i_5_3659 (.A1(n_5_3362), .A2(n_5_2179), .ZN(n_5_3358));
   INV_X1 i_5_3660 (.A(n_5_2234), .ZN(n_5_3361));
   INV_X1 i_5_3661 (.A(n_5_2233), .ZN(n_5_3362));
   INV_X1 i_5_3662 (.A(n_5_2180), .ZN(n_5_3363));
   INV_X1 i_5_3663 (.A(n_5_2179), .ZN(n_5_3368));
   OAI22_X1 i_5_3664 (.A1(n_5_2234), .A2(n_5_3363), .B1(n_5_2233), .B2(n_5_3368), 
      .ZN(n_5_3369));
   OR2_X1 i_5_3665 (.A1(n_5_3418), .A2(m[6]), .ZN(n_5_3370));
   NAND2_X1 i_5_3666 (.A1(n_5_3418), .A2(m[6]), .ZN(n_5_3371));
   XNOR2_X1 i_5_2029 (.A(n_5_3418), .B(m[6]), .ZN(n_5_3373));
   NAND2_X1 i_5_3668 (.A1(n_5_2206), .A2(n_5_3526), .ZN(n_5_3374));
   NAND2_X1 i_5_3669 (.A1(n_5_2206), .A2(n_5_3526), .ZN(n_5_3375));
   XNOR2_X1 i_5_3670 (.A(n_5_3457), .B(n_5_2170), .ZN(n_5_3376));
   NAND2_X1 i_5_3671 (.A1(n_5_3376), .A2(n_5_3386), .ZN(n_5_3378));
   NAND3_X1 i_5_3470 (.A1(n_5_2156), .A2(n_5_2157), .A3(n_5_2158), .ZN(n_5_3382));
   NAND3_X1 i_5_3673 (.A1(n_5_2156), .A2(n_5_2157), .A3(n_5_2158), .ZN(n_5_3388));
   INV_X1 i_5_3674 (.A(n_5_3388), .ZN(n_5_3390));
   INV_X1 i_5_3675 (.A(n_5_2032), .ZN(n_5_3391));
   NAND2_X1 i_5_3676 (.A1(n_5_3390), .A2(n_5_3391), .ZN(n_5_3394));
   INV_X1 i_5_3677 (.A(n_5_2031), .ZN(n_5_3395));
   NAND2_X1 i_5_3678 (.A1(n_5_3388), .A2(n_5_3395), .ZN(n_5_3396));
   NAND2_X1 i_5_3679 (.A1(n_5_3394), .A2(n_5_3396), .ZN(n_5_3400));
   NAND2_X1 i_5_3680 (.A1(n_5_2154), .A2(n_5_3051), .ZN(n_5_3402));
   XNOR2_X1 i_5_3681 (.A(n_5_3402), .B(n_55), .ZN(n_5_3404));
   XNOR2_X1 i_5_3682 (.A(n_5_3402), .B(m[9]), .ZN(n_5_3405));
   NAND2_X1 i_5_3486 (.A1(n_5_2154), .A2(n_5_3051), .ZN(n_5_3406));
   XNOR2_X1 i_5_3684 (.A(n_5_2178), .B(n_5_2225), .ZN(n_5_3407));
   NAND2_X1 i_5_3685 (.A1(n_5_3407), .A2(n_5_3386), .ZN(n_5_3408));
   INV_X1 i_5_3686 (.A(n_5_3150), .ZN(n_5_3409));
   NAND2_X1 i_5_3687 (.A1(n_5_3315), .A2(n_5_3150), .ZN(n_5_3410));
   INV_X1 i_5_3688 (.A(n_5_3410), .ZN(n_5_3411));
   NAND2_X1 i_5_3689 (.A1(n_5_3351), .A2(n_5_3328), .ZN(n_5_3412));
   NAND2_X1 i_5_3690 (.A1(n_5_3351), .A2(n_5_3328), .ZN(n_5_3413));
   INV_X1 i_5_3691 (.A(n_5_3413), .ZN(n_5_3414));
   NAND2_X1 i_5_3692 (.A1(n_5_1212), .A2(n_5_3044), .ZN(n_5_3415));
   INV_X1 i_5_3693 (.A(n_5_3415), .ZN(n_5_3416));
   NAND3_X1 i_5_3694 (.A1(n_5_3378), .A2(n_5_3132), .A3(n_5_3416), .ZN(n_5_3417));
   NAND3_X1 i_5_2055 (.A1(n_5_1213), .A2(n_5_2986), .A3(n_5_2116), .ZN(n_5_3418));
   INV_X1 i_5_3696 (.A(n_5_3185), .ZN(n_5_3419));
   NAND2_X1 i_5_3697 (.A1(n_5_2116), .A2(n_5_3419), .ZN(n_5_3420));
   INV_X1 i_5_3698 (.A(n_5_3420), .ZN(n_5_3421));
   OR3_X1 i_5_3699 (.A1(n_5_3409), .A2(n_5_3424), .A3(n_5_3425), .ZN(n_5_3422));
   INV_X1 i_5_3700 (.A(n_5_3426), .ZN(n_5_3423));
   NOR2_X1 i_5_3701 (.A1(n_5_3063), .A2(n_5_2568), .ZN(n_5_3424));
   NAND2_X1 i_5_3702 (.A1(n_5_1211), .A2(m[0]), .ZN(n_5_3425));
   OAI21_X1 i_5_3703 (.A(n_5_1074), .B1(n_5_3409), .B2(n_5_3057), .ZN(n_5_3426));
   NAND2_X1 i_5_3704 (.A1(n_5_1211), .A2(m[0]), .ZN(n_5_3427));
   INV_X1 i_5_3705 (.A(n_5_3427), .ZN(n_5_3428));
   NAND2_X1 i_5_3706 (.A1(n_5_3063), .A2(n_5_3428), .ZN(n_5_3429));
   NAND2_X1 i_5_3707 (.A1(n_5_2568), .A2(m[0]), .ZN(n_5_3430));
   INV_X1 i_5_3708 (.A(n_5_3430), .ZN(n_5_3431));
   NAND2_X1 i_5_3709 (.A1(n_5_1211), .A2(n_5_3431), .ZN(n_5_3432));
   NAND3_X1 i_5_3710 (.A1(n_5_3057), .A2(n_5_3429), .A3(n_5_3432), .ZN(n_5_3433));
   INV_X1 i_5_3711 (.A(n_5_3433), .ZN(n_5_3434));
   OAI21_X1 i_5_3712 (.A(n_5_1074), .B1(n_5_3434), .B2(n_5_3409), .ZN(n_5_3435));
   INV_X1 i_5_3713 (.A(n_5_3400), .ZN(n_5_3436));
   NAND3_X1 i_5_3714 (.A1(n_5_966), .A2(n_5_1007), .A3(n_5_976), .ZN(n_5_3437));
   NAND2_X1 i_5_3715 (.A1(n_5_982), .A2(n_5_3437), .ZN(n_5_3438));
   NAND3_X1 i_5_3716 (.A1(n_5_966), .A2(n_5_1007), .A3(n_5_976), .ZN(n_5_3439));
   XNOR2_X1 i_5_3717 (.A(n_5_3567), .B(n_5_3027), .ZN(n_5_3440));
   XNOR2_X1 i_5_3718 (.A(n_5_1734), .B(n_5_1778), .ZN(n_5_3441));
   NAND2_X1 i_5_3488 (.A1(n_5_3441), .A2(n_5_3386), .ZN(n_5_3442));
   OAI21_X1 i_5_3720 (.A(n_5_1460), .B1(n_5_3191), .B2(m[13]), .ZN(n_5_4086));
   INV_X1 i_5_3721 (.A(n_5_3375), .ZN(n_5_4087));
   INV_X1 i_5_3722 (.A(m[13]), .ZN(n_5_3443));
   NAND2_X1 i_5_3723 (.A1(n_5_4085), .A2(n_5_3443), .ZN(n_5_3444));
   OAI21_X1 i_5_3724 (.A(n_5_1458), .B1(n_5_3191), .B2(n_5_3444), .ZN(n_5_3445));
   INV_X1 i_5_3725 (.A(n_5_1460), .ZN(n_5_3446));
   AOI21_X1 i_5_3726 (.A(n_5_3445), .B1(n_5_3446), .B2(n_5_4085), .ZN(n_5_3447));
   INV_X1 i_5_3727 (.A(n_5_4085), .ZN(n_5_3448));
   OAI21_X1 i_5_3728 (.A(n_5_3447), .B1(n_5_3375), .B2(n_5_3448), .ZN(n_5_3449));
   NAND2_X1 i_5_3729 (.A1(n_5_3291), .A2(n_60), .ZN(n_5_3450));
   NAND2_X1 i_5_3510 (.A1(n_5_3291), .A2(n_60), .ZN(n_5_3451));
   INV_X1 i_5_3519 (.A(n_5_3451), .ZN(n_5_3452));
   NAND3_X1 i_5_3732 (.A1(n_5_1437), .A2(n_5_1438), .A3(n_5_1439), .ZN(n_5_3453));
   NAND2_X1 i_5_3733 (.A1(n_5_3453), .A2(m[5]), .ZN(n_5_3454));
   NAND3_X1 i_5_3734 (.A1(n_5_3018), .A2(n_5_1787), .A3(n_5_1790), .ZN(n_5_3455));
   NAND2_X1 i_5_3735 (.A1(n_5_1719), .A2(n_58), .ZN(n_5_3456));
   NAND2_X1 i_5_3736 (.A1(n_5_3455), .A2(n_5_3456), .ZN(n_5_3457));
   XNOR2_X1 i_5_3737 (.A(n_5_1286), .B(n_5_1717), .ZN(n_5_3458));
   NAND2_X1 i_5_3738 (.A1(n_5_3458), .A2(n_5_3386), .ZN(n_5_3459));
   NAND2_X1 i_5_3739 (.A1(n_5_3461), .A2(m[4]), .ZN(n_5_3460));
   NAND3_X1 i_5_3740 (.A1(n_5_3462), .A2(n_5_3463), .A3(n_5_1212), .ZN(n_5_3461));
   NAND2_X1 i_5_3741 (.A1(n_5_3237), .A2(n_5_3385), .ZN(n_5_3462));
   NAND2_X1 i_5_3742 (.A1(n_5_3227), .A2(n_5_3386), .ZN(n_5_3463));
   NAND2_X1 i_5_3743 (.A1(n_5_3385), .A2(m[4]), .ZN(n_5_3464));
   INV_X1 i_5_3744 (.A(n_5_3464), .ZN(n_5_3465));
   NAND2_X1 i_5_3745 (.A1(n_5_3237), .A2(n_5_3465), .ZN(n_5_3466));
   NAND2_X1 i_5_3746 (.A1(n_5_3386), .A2(m[4]), .ZN(n_5_3467));
   INV_X1 i_5_3747 (.A(n_5_3467), .ZN(n_5_3468));
   NAND2_X1 i_5_3748 (.A1(n_5_3227), .A2(n_5_3468), .ZN(n_5_3469));
   INV_X1 i_5_3749 (.A(n_5_1212), .ZN(n_5_3470));
   NAND2_X1 i_5_3750 (.A1(n_5_3470), .A2(m[4]), .ZN(n_5_3471));
   NAND3_X1 i_5_3751 (.A1(n_5_3466), .A2(n_5_3469), .A3(n_5_3471), .ZN(n_5_3472));
   INV_X1 i_5_2020 (.A(n_5_1391), .ZN(n_5_3473));
   NAND2_X1 i_5_3753 (.A1(n_5_1143), .A2(n_5_3371), .ZN(n_5_3474));
   NAND2_X1 i_5_3754 (.A1(n_5_3474), .A2(n_5_3370), .ZN(n_5_3475));
   NAND2_X1 i_5_3755 (.A1(n_5_1143), .A2(n_5_3371), .ZN(n_5_3476));
   OAI211_X1 i_5_3756 (.A(n_5_3176), .B(n_5_3177), .C1(n_5_3175), .C2(n_5_3183), 
      .ZN(n_5_3477));
   OAI211_X1 i_5_3757 (.A(n_5_3176), .B(n_5_3177), .C1(n_5_3175), .C2(n_5_3183), 
      .ZN(n_5_3478));
   INV_X1 i_5_3758 (.A(m[11]), .ZN(n_5_3479));
   NAND2_X1 i_5_3759 (.A1(n_5_4067), .A2(n_5_3479), .ZN(n_5_3480));
   INV_X1 i_5_3760 (.A(n_5_3480), .ZN(n_5_3481));
   NAND2_X1 i_5_3761 (.A1(n_5_4464), .A2(n_5_3481), .ZN(n_5_3482));
   INV_X1 i_5_3762 (.A(n_5_3482), .ZN(n_5_3483));
   NAND2_X1 i_5_3763 (.A1(n_5_3483), .A2(n_5_4463), .ZN(n_5_3484));
   NAND2_X1 i_5_3764 (.A1(n_5_3478), .A2(n_5_3484), .ZN(n_5_3485));
   XNOR2_X1 i_5_3765 (.A(n_5_3190), .B(n_5_3182), .ZN(n_5_3486));
   XNOR2_X1 i_5_3766 (.A(n_5_3182), .B(n_5_3190), .ZN(n_5_3487));
   NAND2_X1 i_5_3532 (.A1(n_5_3487), .A2(n_5_3385), .ZN(n_5_3488));
   NAND2_X1 i_5_3768 (.A1(n_5_3180), .A2(n_5_3181), .ZN(n_5_3489));
   INV_X1 i_5_2062 (.A(n_5_3489), .ZN(n_5_3490));
   INV_X1 i_5_3770 (.A(m[6]), .ZN(n_5_3491));
   NAND2_X1 i_5_3771 (.A1(n_5_4653), .A2(n_5_3491), .ZN(n_5_3492));
   INV_X1 i_5_3772 (.A(n_5_3492), .ZN(n_5_3493));
   NAND3_X1 i_5_3773 (.A1(n_5_4659), .A2(n_5_4658), .A3(n_5_3493), .ZN(n_5_3494));
   NAND2_X1 i_5_3774 (.A1(n_5_3138), .A2(n_5_3136), .ZN(n_5_3495));
   INV_X1 i_5_3775 (.A(n_5_420), .ZN(n_5_3496));
   AOI21_X1 i_5_3776 (.A(n_5_3496), .B1(n_5_3136), .B2(n_5_3797), .ZN(n_5_3497));
   NAND2_X1 i_5_3777 (.A1(n_5_3495), .A2(n_5_3497), .ZN(n_5_3498));
   XNOR2_X1 i_5_3778 (.A(n_5_4179), .B(n_5_3131), .ZN(n_5_3499));
   NAND2_X1 i_5_846 (.A1(n_5_3499), .A2(n_5_378), .ZN(n_5_4088));
   NAND2_X1 i_5_3780 (.A1(n_5_3596), .A2(n_5_4017), .ZN(n_5_3500));
   INV_X1 i_5_3781 (.A(n_5_3335), .ZN(n_5_3501));
   AOI21_X1 i_5_3782 (.A(n_5_3501), .B1(n_5_3149), .B2(n_5_1006), .ZN(n_5_3502));
   NAND2_X1 i_5_3783 (.A1(n_5_3158), .A2(n_5_3157), .ZN(n_5_3503));
   NAND2_X1 i_5_3784 (.A1(n_5_3503), .A2(n_5_1038), .ZN(n_5_3504));
   NAND2_X1 i_5_3785 (.A1(n_5_3141), .A2(n_5_3124), .ZN(n_5_3505));
   NAND2_X1 i_5_3786 (.A1(m[3]), .A2(n_5_3139), .ZN(n_5_3506));
   NAND2_X1 i_5_3787 (.A1(m[2]), .A2(n_5_3795), .ZN(n_5_3507));
   NAND2_X1 i_5_3788 (.A1(n_5_3124), .A2(n_5_3141), .ZN(n_5_3508));
   NAND2_X1 i_5_3789 (.A1(n_5_3139), .A2(m[3]), .ZN(n_5_3509));
   NAND2_X1 i_5_3790 (.A1(n_5_3795), .A2(m[2]), .ZN(n_5_3510));
   NAND3_X1 i_5_3791 (.A1(n_5_3508), .A2(n_5_3509), .A3(n_5_3510), .ZN(n_5_3511));
   INV_X1 i_5_3792 (.A(n_5_3128), .ZN(n_5_3512));
   NAND2_X1 i_5_2500 (.A1(n_5_4787), .A2(n_5_3512), .ZN(n_5_3513));
   NAND2_X1 i_5_2501 (.A1(n_5_3933), .A2(m[12]), .ZN(n_5_3514));
   NAND2_X1 i_5_3283 (.A1(n_5_3513), .A2(n_5_3514), .ZN(n_5_3515));
   NAND2_X1 i_5_3796 (.A1(n_5_3168), .A2(m[9]), .ZN(n_5_3516));
   NAND2_X1 i_5_3797 (.A1(n_5_3168), .A2(m[9]), .ZN(n_5_3517));
   OR2_X1 i_5_3798 (.A1(n_5_3418), .A2(n_5_3185), .ZN(n_5_3518));
   NAND2_X1 i_5_3799 (.A1(n_5_3737), .A2(n_5_3738), .ZN(n_5_3519));
   OAI21_X1 i_5_3800 (.A(n_5_3519), .B1(n_5_3418), .B2(n_5_3185), .ZN(n_5_3520));
   INV_X1 i_5_3801 (.A(n_5_3143), .ZN(n_5_3521));
   XNOR2_X1 i_5_3802 (.A(n_5_3209), .B(n_5_3521), .ZN(n_5_3522));
   NAND3_X1 i_5_3803 (.A1(n_5_3164), .A2(n_5_3163), .A3(n_5_3162), .ZN(n_5_3523));
   NAND2_X1 i_5_3804 (.A1(n_5_3188), .A2(n_5_3189), .ZN(n_5_3524));
   NAND2_X1 i_5_3805 (.A1(n_5_3173), .A2(n_5_3174), .ZN(n_5_3525));
   NAND2_X1 i_5_3806 (.A1(n_5_3191), .A2(m[13]), .ZN(n_5_3526));
   NAND2_X1 i_5_3807 (.A1(n_5_3173), .A2(n_5_3174), .ZN(n_5_3527));
   NAND2_X1 i_5_3808 (.A1(n_5_3191), .A2(m[13]), .ZN(n_5_3528));
   NAND2_X1 i_5_3809 (.A1(n_5_3527), .A2(n_5_3528), .ZN(n_5_3529));
   NAND2_X1 i_5_3810 (.A1(n_5_3172), .A2(n_5_3170), .ZN(n_5_3530));
   NAND3_X1 i_5_3811 (.A1(n_5_3723), .A2(n_5_3530), .A3(n_5_3171), .ZN(n_5_464));
   NAND2_X1 i_5_3812 (.A1(n_5_3166), .A2(n_5_3167), .ZN(n_5_3532));
   NAND3_X1 i_5_3813 (.A1(n_5_3517), .A2(n_5_3166), .A3(n_5_3167), .ZN(n_5_3533));
   NAND2_X1 i_5_3814 (.A1(n_5_3165), .A2(n_5_3516), .ZN(n_5_3534));
   NAND2_X1 i_5_3815 (.A1(n_5_3533), .A2(n_5_3534), .ZN(n_5_3535));
   NAND2_X1 i_5_3816 (.A1(n_5_3126), .A2(n_5_3494), .ZN(n_5_3536));
   NAND2_X1 i_5_3817 (.A1(n_5_3129), .A2(n_5_3494), .ZN(n_5_3537));
   NAND2_X1 i_5_3818 (.A1(n_5_3536), .A2(n_5_3537), .ZN(n_5_3538));
   XNOR2_X1 i_5_3819 (.A(n_5_3178), .B(n_5_3179), .ZN(n_5_3539));
   NAND2_X1 i_5_3820 (.A1(n_5_3539), .A2(n_5_1452), .ZN(n_5_3540));
   INV_X1 i_5_3821 (.A(n_5_1791), .ZN(n_5_3541));
   NAND2_X1 i_5_3822 (.A1(n_5_3541), .A2(n_5_2866), .ZN(n_5_3542));
   INV_X1 i_5_3823 (.A(n_5_1716), .ZN(n_5_3543));
   INV_X1 i_5_3824 (.A(n_5_3228), .ZN(n_5_3544));
   NAND2_X1 i_5_3825 (.A1(n_5_3543), .A2(n_5_3544), .ZN(n_5_3545));
   OAI21_X1 i_5_3533 (.A(n_5_3542), .B1(n_5_3545), .B2(n_5_1262), .ZN(n_5_3546));
   NAND3_X1 i_5_3827 (.A1(n_5_1825), .A2(n_5_1827), .A3(n_5_1800), .ZN(n_5_3547));
   XNOR2_X1 i_5_3828 (.A(n_5_3547), .B(n_66), .ZN(n_5_3548));
   NOR2_X1 i_5_3829 (.A1(n_5_3547), .A2(n_66), .ZN(n_5_3549));
   NOR2_X1 i_5_3830 (.A1(n_5_3554), .A2(m[5]), .ZN(n_5_3550));
   NAND2_X1 i_5_3831 (.A1(n_5_3554), .A2(m[5]), .ZN(n_5_3551));
   XNOR2_X1 i_5_3832 (.A(n_5_3547), .B(m[5]), .ZN(n_5_3552));
   NOR2_X1 i_5_3833 (.A1(n_5_3547), .A2(n_66), .ZN(n_5_3553));
   NAND3_X1 i_5_3834 (.A1(n_5_1825), .A2(n_5_1827), .A3(n_5_1800), .ZN(n_5_3554));
   XNOR2_X1 i_5_3835 (.A(n_5_916), .B(n_5_797), .ZN(n_5_3555));
   NAND2_X1 i_5_285 (.A1(n_5_3555), .A2(n_5_378), .ZN(n_5_3556));
   INV_X1 i_5_3837 (.A(n_5_3563), .ZN(n_5_3557));
   NAND2_X1 i_5_3838 (.A1(n_5_4162), .A2(n_5_2568), .ZN(n_5_3558));
   NOR2_X1 i_5_3839 (.A1(n_5_4162), .A2(n_5_2568), .ZN(n_5_3559));
   NAND2_X1 i_5_3840 (.A1(n_5_4162), .A2(n_5_2568), .ZN(n_5_3560));
   NAND2_X1 i_5_3841 (.A1(n_5_4162), .A2(m[1]), .ZN(n_5_3561));
   XNOR2_X1 i_5_3842 (.A(n_5_4162), .B(n_5_736), .ZN(n_5_3562));
   NAND3_X1 i_5_3843 (.A1(n_5_606), .A2(n_5_611), .A3(n_5_605), .ZN(n_5_3563));
   NAND3_X1 i_5_3844 (.A1(n_5_1311), .A2(n_5_3017), .A3(n_5_1785), .ZN(n_5_3564));
   NAND2_X1 i_5_3845 (.A1(n_5_1305), .A2(n_5_1338), .ZN(n_5_3565));
   NAND2_X1 i_5_3846 (.A1(n_5_1784), .A2(n_66), .ZN(n_5_3566));
   NAND3_X1 i_5_3847 (.A1(n_5_3564), .A2(n_5_3565), .A3(n_5_3566), .ZN(n_5_3567));
   NAND2_X1 i_5_3848 (.A1(n_5_3716), .A2(n_5_4017), .ZN(n_5_4656));
   AOI21_X1 i_5_3849 (.A(n_5_653), .B1(n_5_3854), .B2(n_5_1006), .ZN(n_5_4657));
   INV_X1 i_5_2089 (.A(n_5_653), .ZN(n_5_3568));
   NAND3_X1 i_5_2132 (.A1(n_5_3717), .A2(n_5_4588), .A3(n_5_3568), .ZN(n_5_3569));
   NAND3_X1 i_5_3852 (.A1(n_5_2986), .A2(n_5_1213), .A3(n_5_3421), .ZN(n_5_3570));
   INV_X1 i_5_3853 (.A(n_5_3041), .ZN(n_5_3571));
   NAND3_X1 i_5_3854 (.A1(n_5_2986), .A2(n_5_1213), .A3(n_5_3421), .ZN(n_5_3572));
   NAND2_X1 i_5_3855 (.A1(n_5_3571), .A2(n_5_3572), .ZN(n_5_3573));
   NAND3_X1 i_5_3856 (.A1(n_5_1008), .A2(n_5_966), .A3(n_5_976), .ZN(n_5_3574));
   INV_X1 i_5_3857 (.A(n_5_3574), .ZN(n_5_3575));
   INV_X1 i_5_3858 (.A(n_54), .ZN(n_5_3576));
   INV_X1 i_5_3859 (.A(n_5_3704), .ZN(n_5_3577));
   XNOR2_X1 i_5_3860 (.A(n_5_3604), .B(n_5_3703), .ZN(n_5_3578));
   INV_X1 i_5_3861 (.A(n_5_4096), .ZN(n_5_3579));
   AOI21_X1 i_5_3862 (.A(n_5_3749), .B1(n_5_4351), .B2(n_5_3579), .ZN(n_5_3580));
   XNOR2_X1 i_5_3863 (.A(n_5_3626), .B(n_5_3580), .ZN(n_5_3581));
   NOR2_X1 i_5_3864 (.A1(n_5_3401), .A2(n_58), .ZN(n_5_3582));
   INV_X1 i_5_3865 (.A(n_5_3582), .ZN(n_5_3583));
   NAND2_X1 i_5_3866 (.A1(n_5_3401), .A2(n_58), .ZN(n_5_3584));
   INV_X1 i_5_3867 (.A(n_5_3584), .ZN(n_5_3585));
   OAI21_X1 i_5_3868 (.A(n_5_3583), .B1(n_5_3585), .B2(n_5_3629), .ZN(n_5_3586));
   AOI21_X1 i_5_3869 (.A(n_5_3652), .B1(n_5_3586), .B2(n_5_4148), .ZN(n_5_4089));
   AOI21_X1 i_5_3870 (.A(n_5_3611), .B1(n_5_3690), .B2(n_5_3653), .ZN(n_5_3587));
   INV_X1 i_5_3871 (.A(n_5_4139), .ZN(n_5_4090));
   INV_X1 i_5_3872 (.A(n_5_3666), .ZN(n_5_3588));
   OAI21_X1 i_5_3534 (.A(n_5_3665), .B1(n_5_3610), .B2(n_5_3588), .ZN(n_5_4091));
   NOR2_X1 i_5_3874 (.A1(n_5_3377), .A2(n_61), .ZN(n_5_3589));
   INV_X1 i_5_3875 (.A(n_5_3589), .ZN(n_5_4092));
   NAND2_X1 i_5_3876 (.A1(n_5_3377), .A2(n_61), .ZN(n_5_4093));
   OR2_X1 i_5_3877 (.A1(n_5_3399), .A2(n_53), .ZN(n_5_3590));
   NAND2_X1 i_5_3878 (.A1(n_5_3399), .A2(n_53), .ZN(n_5_3591));
   NAND2_X1 i_5_3879 (.A1(n_5_3590), .A2(n_5_3591), .ZN(n_5_3592));
   NAND3_X1 i_5_3880 (.A1(n_5_3605), .A2(n_5_3701), .A3(n_5_4093), .ZN(n_5_3593));
   NAND3_X1 i_5_3881 (.A1(n_5_3592), .A2(n_5_4092), .A3(n_5_3593), .ZN(n_5_3594));
   AOI21_X1 i_5_3882 (.A(n_5_3589), .B1(n_5_4510), .B2(n_5_4093), .ZN(n_5_3595));
   OAI21_X1 i_5_3883 (.A(n_5_3594), .B1(n_5_3592), .B2(n_5_3595), .ZN(n_5_3596));
   XNOR2_X1 i_5_3884 (.A(n_5_3576), .B(n_53), .ZN(n_5_3597));
   NAND2_X1 i_5_3885 (.A1(n_5_3590), .A2(n_5_4093), .ZN(n_5_3598));
   NAND2_X1 i_5_3886 (.A1(n_5_4092), .A2(n_5_3700), .ZN(n_5_3599));
   INV_X1 i_5_3887 (.A(n_5_3634), .ZN(n_5_3600));
   AOI21_X1 i_5_3888 (.A(n_5_3599), .B1(n_5_3600), .B2(n_5_3701), .ZN(n_5_3601));
   INV_X1 i_5_3889 (.A(n_5_3599), .ZN(n_5_3602));
   NAND3_X1 i_5_3890 (.A1(n_5_3701), .A2(n_5_3985), .A3(n_5_3656), .ZN(n_5_3603));
   INV_X1 i_5_3891 (.A(n_5_3749), .ZN(n_5_4094));
   XNOR2_X1 i_5_3892 (.A(n_5_4101), .B(n_59), .ZN(n_5_3604));
   NAND2_X1 i_5_3893 (.A1(n_5_3700), .A2(n_5_3634), .ZN(n_5_3605));
   INV_X1 i_5_3894 (.A(n_5_4108), .ZN(n_5_3606));
   INV_X1 i_5_3895 (.A(n_55), .ZN(n_5_3607));
   NAND2_X1 i_5_3896 (.A1(n_5_3606), .A2(n_5_3607), .ZN(n_5_3608));
   NAND2_X1 i_5_3897 (.A1(n_5_3677), .A2(n_5_3608), .ZN(n_5_3609));
   NAND2_X1 i_5_3898 (.A1(n_5_3609), .A2(n_5_3715), .ZN(n_5_3610));
   NOR2_X1 i_5_3899 (.A1(n_5_4192), .A2(n_5_3185), .ZN(n_5_3611));
   INV_X1 i_5_3900 (.A(n_5_3185), .ZN(n_5_3612));
   NAND2_X1 i_5_3901 (.A1(n_5_3365), .A2(n_5_2568), .ZN(n_5_3613));
   NAND2_X1 i_5_3902 (.A1(n_5_3364), .A2(m[0]), .ZN(n_5_3614));
   NAND2_X1 i_5_3903 (.A1(n_5_2568), .A2(m[0]), .ZN(n_5_3615));
   INV_X1 i_5_3904 (.A(n_5_3615), .ZN(n_5_3616));
   NAND2_X1 i_5_3905 (.A1(n_5_3364), .A2(n_5_3616), .ZN(n_5_3617));
   INV_X1 i_5_3906 (.A(n_5_3617), .ZN(n_5_3618));
   NOR2_X1 i_5_3907 (.A1(n_5_2568), .A2(m[0]), .ZN(n_5_3619));
   INV_X1 i_5_3908 (.A(n_5_3364), .ZN(n_5_3620));
   INV_X1 i_5_3909 (.A(n_5_2568), .ZN(n_5_3621));
   AOI21_X1 i_5_3910 (.A(n_5_3619), .B1(n_5_3620), .B2(n_5_3621), .ZN(n_5_3622));
   NAND2_X1 i_5_3911 (.A1(n_5_3625), .A2(n_5_3684), .ZN(n_5_3623));
   NAND2_X1 i_5_3912 (.A1(n_5_4385), .A2(n_5_3623), .ZN(n_5_3624));
   INV_X1 i_5_3913 (.A(n_5_3804), .ZN(n_5_4095));
   NOR2_X1 i_5_3914 (.A1(n_5_3381), .A2(n_65), .ZN(n_5_3625));
   XNOR2_X1 i_5_3915 (.A(n_5_3381), .B(n_65), .ZN(n_5_3626));
   NAND2_X1 i_5_3916 (.A1(n_5_4194), .A2(n_5_3612), .ZN(n_5_3627));
   INV_X1 i_5_3917 (.A(n_5_3627), .ZN(n_5_3628));
   OAI21_X1 i_5_3918 (.A(n_5_3684), .B1(n_5_3625), .B2(n_5_3683), .ZN(n_5_3629));
   INV_X1 i_5_3919 (.A(n_5_3583), .ZN(n_5_3630));
   NAND2_X1 i_5_3920 (.A1(n_5_3365), .A2(n_5_3622), .ZN(n_5_3631));
   INV_X1 i_5_3921 (.A(n_5_3618), .ZN(n_5_3633));
   NAND2_X1 i_5_3922 (.A1(n_5_3631), .A2(n_5_3633), .ZN(n_5_4096));
   NAND2_X1 i_5_3923 (.A1(n_5_3656), .A2(n_5_3985), .ZN(n_5_3634));
   NAND2_X1 i_5_3924 (.A1(n_5_3372), .A2(n_69), .ZN(n_5_3635));
   NOR2_X1 i_5_3925 (.A1(n_5_3372), .A2(n_69), .ZN(n_5_3636));
   XNOR2_X1 i_5_3926 (.A(n_5_3372), .B(n_69), .ZN(n_5_3637));
   AOI21_X1 i_5_3927 (.A(n_5_4353), .B1(n_5_4094), .B2(n_5_4096), .ZN(n_5_3638));
   OAI21_X1 i_5_3928 (.A(n_5_3684), .B1(n_5_3638), .B2(n_5_3625), .ZN(n_5_3640));
   INV_X1 i_5_3929 (.A(n_5_4481), .ZN(n_5_3641));
   INV_X1 i_5_3930 (.A(n_5_3714), .ZN(n_5_3642));
   OAI21_X1 i_5_3931 (.A(n_5_4139), .B1(n_5_3678), .B2(n_5_3804), .ZN(n_5_3643));
   NAND2_X1 i_5_3932 (.A1(n_5_3636), .A2(n_5_3635), .ZN(n_5_3644));
   INV_X1 i_5_3933 (.A(n_5_3635), .ZN(n_5_3645));
   INV_X1 i_5_3934 (.A(n_5_4155), .ZN(n_5_3646));
   INV_X1 i_5_3935 (.A(n_73), .ZN(n_5_3647));
   NAND2_X1 i_5_3936 (.A1(n_5_3646), .A2(n_5_3647), .ZN(n_5_3648));
   NAND2_X1 i_5_3937 (.A1(n_5_3648), .A2(n_5_3643), .ZN(n_5_3649));
   INV_X1 i_5_3938 (.A(n_5_3649), .ZN(n_5_3650));
   INV_X1 i_5_3939 (.A(n_5_4154), .ZN(n_5_3651));
   NOR2_X1 i_5_3940 (.A1(n_5_4150), .A2(n_66), .ZN(n_5_3652));
   NAND2_X1 i_5_3941 (.A1(n_5_4192), .A2(n_5_3185), .ZN(n_5_3653));
   NAND2_X1 i_5_3942 (.A1(n_5_4194), .A2(n_5_3612), .ZN(n_5_3654));
   NAND2_X1 i_5_3943 (.A1(n_5_4192), .A2(n_5_3185), .ZN(n_5_3655));
   NAND2_X1 i_5_3944 (.A1(n_5_3654), .A2(n_5_3655), .ZN(n_5_4097));
   NAND2_X1 i_5_709 (.A1(n_5_3680), .A2(n_5_3675), .ZN(n_5_3656));
   NOR2_X1 i_5_3946 (.A1(n_76), .A2(n_75), .ZN(n_5_3657));
   INV_X1 i_5_3947 (.A(n_5_3983), .ZN(n_5_3658));
   INV_X1 i_5_3948 (.A(n_75), .ZN(n_5_3659));
   NAND2_X1 i_5_3949 (.A1(n_76), .A2(n_75), .ZN(n_5_3660));
   INV_X1 i_5_3950 (.A(n_5_3660), .ZN(n_5_3661));
   NAND2_X1 i_5_3951 (.A1(n_5_3983), .A2(n_5_3661), .ZN(n_5_3662));
   OAI21_X1 i_5_3952 (.A(n_5_3635), .B1(n_5_3668), .B2(n_5_3636), .ZN(n_5_3663));
   XNOR2_X1 i_5_3953 (.A(n_5_4138), .B(n_5_3663), .ZN(n_5_3664));
   OAI21_X1 i_5_3954 (.A(n_5_3635), .B1(n_5_3668), .B2(n_5_3636), .ZN(n_5_4098));
   INV_X1 i_5_3955 (.A(n_5_3667), .ZN(n_5_3665));
   NAND2_X1 i_5_3956 (.A1(n_5_4155), .A2(n_73), .ZN(n_5_3666));
   NOR2_X1 i_5_3957 (.A1(n_5_4155), .A2(n_73), .ZN(n_5_3667));
   NAND2_X1 i_5_3958 (.A1(n_5_3693), .A2(n_5_3694), .ZN(n_5_3668));
   INV_X1 i_5_3959 (.A(n_5_3614), .ZN(n_5_3669));
   XNOR2_X1 i_5_3960 (.A(n_5_3613), .B(n_5_3669), .ZN(n_5_3670));
   INV_X1 i_5_3961 (.A(n_5_3577), .ZN(n_5_3671));
   OAI22_X1 i_5_3962 (.A1(n_5_3670), .A2(n_5_3671), .B1(n_5_3577), .B2(n_5_3614), 
      .ZN(n_5_3672));
   NAND2_X1 i_5_3963 (.A1(n_5_3650), .A2(n_5_3642), .ZN(n_5_3673));
   AOI21_X1 i_5_3964 (.A(n_5_3651), .B1(n_5_3641), .B2(n_5_3648), .ZN(n_5_3674));
   NAND2_X1 i_5_3965 (.A1(n_5_3673), .A2(n_5_3674), .ZN(n_5_3675));
   OAI21_X1 i_5_3966 (.A(n_5_3644), .B1(n_5_3695), .B2(n_5_3645), .ZN(n_5_3676));
   OAI21_X1 i_5_3967 (.A(n_5_4139), .B1(n_5_3804), .B2(n_5_3676), .ZN(n_5_3677));
   OAI21_X1 i_5_3968 (.A(n_5_3644), .B1(n_5_3695), .B2(n_5_3645), .ZN(n_5_3678));
   OAI211_X1 i_5_3969 (.A(n_5_3680), .B(n_5_3675), .C1(n_5_678), .C2(n_75), 
      .ZN(n_5_3679));
   NAND2_X1 i_5_3970 (.A1(n_5_3679), .A2(n_5_3713), .ZN(n_5_4099));
   OR2_X1 i_5_3971 (.A1(n_5_3983), .A2(n_76), .ZN(n_5_3680));
   AOI21_X1 i_5_3973 (.A(n_5_4353), .B1(n_5_4094), .B2(n_5_4096), .ZN(n_5_3683));
   NAND2_X1 i_5_3974 (.A1(n_5_3381), .A2(n_65), .ZN(n_5_3684));
   NAND2_X1 i_5_3975 (.A1(n_5_3381), .A2(n_65), .ZN(n_5_3685));
   OAI21_X1 i_5_3976 (.A(n_5_3584), .B1(n_5_3624), .B2(n_5_3582), .ZN(n_5_3686));
   NAND2_X1 i_5_3977 (.A1(n_5_3652), .A2(n_5_4148), .ZN(n_5_3687));
   NOR2_X1 i_5_3978 (.A1(n_5_3582), .A2(n_5_3624), .ZN(n_5_3688));
   NAND2_X1 i_5_3979 (.A1(n_5_4148), .A2(n_5_3584), .ZN(n_5_3689));
   OAI21_X1 i_5_3980 (.A(n_5_3687), .B1(n_5_3688), .B2(n_5_3689), .ZN(n_5_3690));
   NAND2_X1 i_5_3981 (.A1(n_5_3591), .A2(n_5_3597), .ZN(n_5_3691));
   INV_X1 i_5_3982 (.A(n_5_3691), .ZN(n_5_3692));
   NAND2_X1 i_5_3983 (.A1(n_5_3628), .A2(n_5_3653), .ZN(n_5_3693));
   NAND2_X1 i_5_3984 (.A1(n_5_3690), .A2(n_5_3653), .ZN(n_5_3694));
   OAI21_X1 i_5_3985 (.A(n_5_3653), .B1(n_5_3628), .B2(n_5_3690), .ZN(n_5_3695));
   NAND2_X1 i_5_3986 (.A1(n_5_3598), .A2(n_5_3591), .ZN(n_5_3696));
   NAND2_X1 i_5_3987 (.A1(n_5_3591), .A2(n_5_3603), .ZN(n_5_3697));
   INV_X1 i_5_3988 (.A(n_5_3697), .ZN(n_5_3698));
   NAND2_X1 i_5_3989 (.A1(n_5_3602), .A2(n_5_3698), .ZN(n_5_3699));
   OR2_X1 i_5_3990 (.A1(n_5_678), .A2(n_75), .ZN(n_5_3700));
   NAND2_X1 i_5_3991 (.A1(n_5_678), .A2(n_75), .ZN(n_5_3701));
   NOR2_X1 i_5_3992 (.A1(n_5_3365), .A2(n_5_2568), .ZN(n_5_3702));
   AOI21_X1 i_5_3993 (.A(n_5_3702), .B1(n_5_3613), .B2(n_5_3614), .ZN(n_5_3703));
   NOR2_X1 i_5_3994 (.A1(n_5_3365), .A2(n_5_2568), .ZN(n_5_3704));
   XNOR2_X1 i_5_719 (.A(n_5_678), .B(n_75), .ZN(n_5_476));
   INV_X1 i_5_729 (.A(n_5_3656), .ZN(n_5_486));
   XNOR2_X1 i_5_737 (.A(n_5_3985), .B(n_75), .ZN(n_5_497));
   NAND2_X1 i_5_4001 (.A1(n_5_3685), .A2(n_5_4351), .ZN(n_5_4100));
   AOI21_X1 i_5_4002 (.A(n_5_3657), .B1(n_5_3658), .B2(n_5_3659), .ZN(n_5_3711));
   INV_X1 i_5_4003 (.A(n_5_3662), .ZN(n_5_3712));
   OAI21_X1 i_5_4004 (.A(n_5_3711), .B1(n_5_678), .B2(n_5_3712), .ZN(n_5_3713));
   NOR2_X1 i_5_4005 (.A1(n_5_4108), .A2(n_55), .ZN(n_5_3714));
   NAND2_X1 i_5_4006 (.A1(n_5_4108), .A2(n_55), .ZN(n_5_3715));
   XNOR2_X1 i_5_4007 (.A(n_5_3900), .B(n_5_4573), .ZN(n_5_3716));
   NAND2_X1 i_5_2160 (.A1(n_5_3896), .A2(n_5_4017), .ZN(n_5_3717));
   NAND2_X1 i_5_4009 (.A1(n_5_4167), .A2(n_5_3340), .ZN(n_5_3718));
   INV_X1 i_5_695 (.A(n_5_3332), .ZN(n_5_3719));
   INV_X1 i_5_699 (.A(n_5_3332), .ZN(n_5_3720));
   INV_X1 i_5_4012 (.A(n_5_1452), .ZN(n_5_3721));
   AOI21_X1 i_5_4013 (.A(n_5_3721), .B1(n_5_4455), .B2(n_5_3403), .ZN(n_5_3722));
   NAND2_X1 i_5_4014 (.A1(n_5_4456), .A2(n_5_3722), .ZN(n_5_3723));
   NAND2_X1 i_5_4015 (.A1(n_5_3833), .A2(n_5_4017), .ZN(n_5_3724));
   INV_X1 i_5_4016 (.A(n_5_3335), .ZN(n_5_3725));
   AOI21_X1 i_5_4017 (.A(n_5_3725), .B1(n_5_3522), .B2(n_5_3333), .ZN(n_5_3726));
   NAND2_X1 i_5_4018 (.A1(n_5_3724), .A2(n_5_3726), .ZN(n_5_3727));
   XNOR2_X1 i_5_4019 (.A(n_5_3848), .B(n_5_3677), .ZN(n_5_3728));
   NAND2_X1 i_5_4020 (.A1(n_5_3728), .A2(n_5_4017), .ZN(n_5_3729));
   NAND2_X1 i_5_4021 (.A1(n_5_3392), .A2(n_5_4069), .ZN(n_5_3730));
   NAND2_X1 i_5_4022 (.A1(n_5_3393), .A2(n_5_4068), .ZN(n_5_3731));
   INV_X1 i_5_4023 (.A(n_5_3389), .ZN(n_5_3732));
   NAND3_X1 i_5_2177 (.A1(n_5_3730), .A2(n_5_3731), .A3(n_5_3732), .ZN(n_5_3733));
   NAND2_X1 i_5_4025 (.A1(n_5_3350), .A2(n_5_4116), .ZN(n_5_3734));
   OAI21_X1 i_5_700 (.A(n_5_4115), .B1(n_5_4323), .B2(n_5_3352), .ZN(n_5_3735));
   NAND2_X1 i_5_4027 (.A1(n_5_3380), .A2(n_5_3397), .ZN(n_5_3737));
   NAND2_X1 i_5_4028 (.A1(n_5_3398), .A2(n_65), .ZN(n_5_3738));
   NAND2_X1 i_5_4029 (.A1(n_5_3397), .A2(n_5_3380), .ZN(n_5_3739));
   NAND2_X1 i_5_4030 (.A1(n_5_3398), .A2(n_65), .ZN(n_5_3740));
   NAND2_X1 i_5_4031 (.A1(n_5_3739), .A2(n_5_3740), .ZN(n_5_3741));
   NAND2_X1 i_5_4032 (.A1(n_5_3387), .A2(n_5_3385), .ZN(n_5_3742));
   NAND2_X1 i_5_4033 (.A1(n_5_3440), .A2(n_5_3386), .ZN(n_5_3743));
   NAND2_X1 i_5_4034 (.A1(n_5_3387), .A2(n_5_3385), .ZN(n_5_3744));
   NAND2_X1 i_5_4035 (.A1(n_5_3440), .A2(n_5_3386), .ZN(n_5_3745));
   NAND3_X1 i_5_4036 (.A1(n_5_3744), .A2(n_5_3745), .A3(n_5_3384), .ZN(n_5_3746));
   XNOR2_X1 i_5_4037 (.A(n_5_3357), .B(n_5_3360), .ZN(n_5_3747));
   NAND2_X1 i_5_701 (.A1(n_5_3747), .A2(n_5_3345), .ZN(n_5_4658));
   NAND3_X1 i_5_4039 (.A1(n_5_3366), .A2(n_5_3383), .A3(n_5_3367), .ZN(n_5_3748));
   NOR2_X1 i_5_4040 (.A1(n_5_3748), .A2(n_59), .ZN(n_5_3749));
   XNOR2_X1 i_5_4041 (.A(n_5_4101), .B(m[2]), .ZN(n_5_3750));
   NOR2_X1 i_5_4042 (.A1(n_5_3748), .A2(m[2]), .ZN(n_5_3751));
   NAND3_X1 i_5_4043 (.A1(n_5_3366), .A2(n_5_3383), .A3(n_5_3367), .ZN(n_5_4101));
   XNOR2_X1 i_5_4044 (.A(n_5_3587), .B(n_5_3637), .ZN(n_5_3752));
   NAND2_X1 i_5_711 (.A1(n_5_3752), .A2(n_5_4017), .ZN(n_5_4659));
   NAND3_X1 i_5_4046 (.A1(n_5_1020), .A2(n_5_1019), .A3(n_5_1021), .ZN(n_5_3753));
   NAND2_X1 i_5_4047 (.A1(n_5_3753), .A2(n_5_3359), .ZN(n_5_3754));
   XNOR2_X1 i_5_4048 (.A(n_5_4237), .B(n_5_3347), .ZN(n_5_3755));
   NAND2_X1 i_5_850 (.A1(n_5_3755), .A2(n_5_420), .ZN(n_5_4102));
   XNOR2_X1 i_5_4050 (.A(n_5_3355), .B(n_5_3356), .ZN(n_5_3756));
   NAND2_X1 i_5_4051 (.A1(n_5_3756), .A2(n_5_3338), .ZN(n_5_3757));
   XNOR2_X1 i_5_4052 (.A(n_5_3341), .B(n_5_3339), .ZN(n_5_3758));
   NAND2_X1 i_5_4053 (.A1(n_5_3758), .A2(n_5_378), .ZN(n_5_4103));
   XNOR2_X1 i_5_4054 (.A(n_5_2699), .B(n_5_3337), .ZN(n_5_3759));
   NAND2_X1 i_5_716 (.A1(n_5_3759), .A2(n_5_635), .ZN(n_5_3760));
   NAND3_X1 i_5_4056 (.A1(n_5_3343), .A2(n_5_4175), .A3(n_5_4238), .ZN(n_5_3761));
   NAND2_X1 i_5_4057 (.A1(m[4]), .A2(n_5_3919), .ZN(n_5_3762));
   NAND3_X1 i_5_4058 (.A1(n_5_4238), .A2(n_5_3343), .A3(n_5_4175), .ZN(n_5_3763));
   NAND2_X1 i_5_4059 (.A1(n_5_3919), .A2(m[4]), .ZN(n_5_3764));
   XNOR2_X1 i_5_4060 (.A(n_5_3741), .B(n_5_3379), .ZN(n_5_3765));
   NAND2_X1 i_5_4061 (.A1(n_5_3765), .A2(n_5_1038), .ZN(n_5_3766));
   NAND3_X1 i_5_732 (.A1(n_5_4659), .A2(n_5_4658), .A3(n_5_4653), .ZN(n_5_3767));
   XNOR2_X1 i_5_4063 (.A(n_5_3767), .B(n_5_841), .ZN(n_5_3768));
   XNOR2_X1 i_5_735 (.A(n_5_3767), .B(n_5_841), .ZN(n_5_3769));
   NAND2_X1 i_5_4065 (.A1(m[6]), .A2(n_5_3767), .ZN(n_5_3770));
   XNOR2_X1 i_5_4066 (.A(n_5_3767), .B(m[6]), .ZN(n_5_873));
   XNOR2_X1 i_5_4067 (.A(n_5_3436), .B(n_5_1142), .ZN(n_5_3772));
   NAND2_X1 i_5_2179 (.A1(n_5_3772), .A2(n_5_1036), .ZN(n_5_3773));
   XNOR2_X1 i_5_4069 (.A(n_5_4097), .B(n_5_4089), .ZN(n_5_3774));
   NAND2_X1 i_5_741 (.A1(n_5_3774), .A2(n_5_4017), .ZN(n_5_3775));
   INV_X1 i_5_4071 (.A(n_5_3795), .ZN(n_5_3776));
   INV_X1 i_5_4072 (.A(n_5_674), .ZN(n_5_3777));
   NOR2_X1 i_5_4073 (.A1(n_5_3795), .A2(n_5_3777), .ZN(n_5_3778));
   NAND2_X1 i_5_759 (.A1(n_5_3919), .A2(n_58), .ZN(n_5_4104));
   NOR2_X1 i_5_4075 (.A1(n_5_858), .A2(n_5_866), .ZN(n_5_3779));
   NAND2_X1 i_5_4076 (.A1(n_5_4042), .A2(n_5_4044), .ZN(n_5_3780));
   NAND2_X1 i_5_4077 (.A1(n_5_3919), .A2(n_58), .ZN(n_5_3781));
   AOI21_X1 i_5_4078 (.A(n_5_3779), .B1(n_5_3780), .B2(n_5_3781), .ZN(n_5_3782));
   NAND2_X1 i_5_4079 (.A1(n_5_3500), .A2(n_5_3502), .ZN(n_5_3783));
   XNOR2_X1 i_5_4080 (.A(m[13]), .B(n_5_3783), .ZN(n_5_3784));
   XNOR2_X1 i_5_4081 (.A(n_5_3783), .B(n_5_751), .ZN(n_5_3785));
   NAND2_X1 i_5_4082 (.A1(n_5_3783), .A2(n_61), .ZN(n_5_3786));
   INV_X1 i_5_4083 (.A(n_5_3783), .ZN(n_5_3787));
   XNOR2_X1 i_5_4084 (.A(n_5_1141), .B(n_5_1130), .ZN(n_5_3788));
   NAND2_X1 i_5_2180 (.A1(n_5_3788), .A2(n_5_1036), .ZN(n_5_3789));
   XNOR2_X1 i_5_4086 (.A(n_5_3035), .B(n_5_1047), .ZN(n_5_3790));
   NAND2_X1 i_5_4087 (.A1(n_5_3790), .A2(n_5_1038), .ZN(n_5_3791));
   NOR2_X1 i_5_2300 (.A1(n_5_3793), .A2(n_69), .ZN(n_5_3792));
   NAND3_X1 i_5_4089 (.A1(n_5_4004), .A2(n_5_4014), .A3(n_5_4016), .ZN(n_5_3793));
   NAND2_X1 i_5_909 (.A1(n_5_3757), .A2(n_5_652), .ZN(n_5_3794));
   NAND2_X1 i_5_4091 (.A1(n_5_3757), .A2(n_5_652), .ZN(n_5_3795));
   NAND2_X1 i_5_1012 (.A1(n_5_3794), .A2(n_59), .ZN(n_5_3796));
   NOR2_X1 i_5_1125 (.A1(n_5_3794), .A2(n_59), .ZN(n_5_3797));
   XNOR2_X1 i_5_4094 (.A(n_5_3794), .B(m[2]), .ZN(n_5_3798));
   XNOR2_X1 i_5_1165 (.A(n_5_907), .B(n_5_866), .ZN(n_5_3799));
   NAND2_X1 i_5_1176 (.A1(n_5_3799), .A2(n_5_420), .ZN(n_5_3865));
   INV_X1 i_5_4097 (.A(n_60), .ZN(n_5_3800));
   NAND2_X1 i_5_4098 (.A1(n_5_1026), .A2(n_5_3800), .ZN(n_5_3801));
   INV_X1 i_5_4099 (.A(n_5_3801), .ZN(n_5_3802));
   NAND3_X1 i_5_4100 (.A1(n_5_1024), .A2(n_5_1025), .A3(n_5_3802), .ZN(n_5_3803));
   INV_X1 i_5_4101 (.A(n_5_3803), .ZN(n_5_3804));
   NAND2_X1 i_5_4102 (.A1(n_5_623), .A2(n_5_621), .ZN(n_5_3805));
   INV_X1 i_5_4103 (.A(n_5_3805), .ZN(n_5_498));
   XNOR2_X1 i_5_4106 (.A(n_5_1751), .B(n_5_1299), .ZN(n_5_3810));
   NOR2_X1 i_5_4107 (.A1(n_5_1284), .A2(n_5_1283), .ZN(n_5_3811));
   NAND2_X1 i_5_4108 (.A1(n_5_3810), .A2(n_5_3811), .ZN(n_5_3812));
   NAND3_X1 i_5_4109 (.A1(n_5_1314), .A2(n_5_1317), .A3(n_5_1315), .ZN(n_5_3813));
   INV_X1 i_5_4110 (.A(n_5_1751), .ZN(n_5_3814));
   XNOR2_X1 i_5_4111 (.A(n_5_3813), .B(n_5_3814), .ZN(n_5_3815));
   OAI21_X1 i_5_4112 (.A(n_5_3812), .B1(n_5_3815), .B2(n_5_3811), .ZN(n_5_3816));
   NAND2_X1 i_5_908 (.A1(n_5_3901), .A2(n_5_4017), .ZN(n_5_3817));
   NAND2_X1 i_5_910 (.A1(n_5_3825), .A2(n_5_640), .ZN(n_5_3818));
   NAND2_X1 i_5_3570 (.A1(n_5_3524), .A2(n_5_3523), .ZN(n_5_3819));
   NOR2_X1 i_5_3601 (.A1(n_5_3115), .A2(n_5_3093), .ZN(n_5_3820));
   NAND2_X1 i_5_3602 (.A1(n_5_3819), .A2(n_5_3820), .ZN(n_5_3821));
   NAND3_X1 i_5_4118 (.A1(n_5_1831), .A2(n_5_1832), .A3(n_5_1799), .ZN(n_5_3822));
   INV_X1 i_5_4119 (.A(m[2]), .ZN(n_5_3823));
   NAND4_X1 i_5_4120 (.A1(n_5_1831), .A2(n_5_1832), .A3(n_5_1799), .A4(n_5_3823), 
      .ZN(n_5_3824));
   XNOR2_X1 i_5_4121 (.A(n_5_1003), .B(n_5_4147), .ZN(n_5_3825));
   XNOR2_X1 i_5_4122 (.A(n_5_4147), .B(n_5_1003), .ZN(n_5_3826));
   NAND2_X1 i_5_4123 (.A1(n_5_3826), .A2(n_5_640), .ZN(n_5_4107));
   NAND2_X1 i_5_4124 (.A1(n_5_3630), .A2(n_5_3640), .ZN(n_5_3827));
   XNOR2_X1 i_5_4125 (.A(n_5_3584), .B(n_5_3640), .ZN(n_5_3828));
   OAI21_X1 i_5_1177 (.A(n_5_3827), .B1(n_5_3828), .B2(n_5_3630), .ZN(n_5_3829));
   INV_X1 i_5_4127 (.A(n_5_3597), .ZN(n_5_3830));
   NAND3_X1 i_5_4128 (.A1(n_5_3699), .A2(n_5_3696), .A3(n_5_3830), .ZN(n_5_3831));
   OAI21_X1 i_5_4129 (.A(n_5_3692), .B1(n_5_3601), .B2(n_5_3598), .ZN(n_5_3832));
   NAND2_X1 i_5_4130 (.A1(n_5_3831), .A2(n_5_3832), .ZN(n_5_3833));
   INV_X1 i_5_4131 (.A(n_63), .ZN(n_5_3834));
   INV_X1 i_5_4132 (.A(n_56), .ZN(n_5_3835));
   NAND2_X1 i_5_4133 (.A1(n_63), .A2(n_56), .ZN(n_5_3836));
   NAND2_X1 i_5_4134 (.A1(n_57), .A2(m[0]), .ZN(n_5_3837));
   NAND2_X1 i_5_4135 (.A1(n_5_3836), .A2(n_5_3837), .ZN(n_5_3838));
   NAND3_X1 i_5_2301 (.A1(n_5_964), .A2(n_5_997), .A3(n_5_959), .ZN(n_5_3842));
   NAND3_X1 i_5_4140 (.A1(n_5_964), .A2(n_5_997), .A3(n_5_959), .ZN(n_5_3843));
   OAI21_X1 i_5_3607 (.A(n_5_4137), .B1(n_5_3843), .B2(n_5_970), .ZN(n_5_3844));
   OAI21_X1 i_5_2303 (.A(n_5_4137), .B1(n_5_3842), .B2(n_5_970), .ZN(n_5_3845));
   XNOR2_X1 i_5_4143 (.A(n_5_3843), .B(n_5_4136), .ZN(n_5_3846));
   NAND3_X1 i_5_2483 (.A1(n_5_3773), .A2(n_5_1027), .A3(n_5_1028), .ZN(n_5_3847));
   XNOR2_X1 i_5_4145 (.A(n_5_3847), .B(n_55), .ZN(n_5_3848));
   NOR2_X1 i_5_2484 (.A1(n_5_3847), .A2(m[9]), .ZN(n_5_3849));
   XNOR2_X1 i_5_4147 (.A(n_5_3847), .B(n_5_992), .ZN(n_5_3850));
   NAND3_X1 i_5_2497 (.A1(n_5_3773), .A2(n_5_1027), .A3(n_5_1028), .ZN(n_5_4108));
   NAND2_X1 i_5_4149 (.A1(n_5_1705), .A2(n_5_1735), .ZN(n_5_3851));
   NAND3_X1 i_5_4150 (.A1(n_5_1736), .A2(n_5_1754), .A3(n_5_1737), .ZN(n_5_3852));
   NAND2_X1 i_5_4151 (.A1(n_5_3851), .A2(n_5_3852), .ZN(n_5_3853));
   XNOR2_X1 i_5_4152 (.A(n_5_3870), .B(n_5_3864), .ZN(n_5_3854));
   XNOR2_X1 i_5_4153 (.A(n_5_4155), .B(m[10]), .ZN(n_5_3870));
   NAND2_X1 i_5_4154 (.A1(n_5_3500), .A2(n_5_3502), .ZN(n_5_3884));
   NAND3_X1 i_5_4155 (.A1(n_5_760), .A2(n_5_757), .A3(n_5_756), .ZN(n_5_3885));
   AOI22_X1 i_5_4156 (.A1(n_5_4787), .A2(n_5_762), .B1(n_5_3500), .B2(n_5_3502), 
      .ZN(n_5_3892));
   NAND2_X1 i_5_4157 (.A1(n_5_3885), .A2(n_5_3892), .ZN(n_5_3894));
   XNOR2_X1 i_5_2499 (.A(n_5_4573), .B(n_5_4153), .ZN(n_5_3896));
   XNOR2_X1 i_5_4159 (.A(n_5_4155), .B(n_73), .ZN(n_5_3900));
   XNOR2_X1 i_5_4160 (.A(n_5_4149), .B(n_5_3686), .ZN(n_5_3901));
   XNOR2_X1 i_5_4161 (.A(n_5_3686), .B(n_5_4149), .ZN(n_5_3902));
   NAND2_X1 i_5_4162 (.A1(n_5_3902), .A2(n_5_4017), .ZN(n_5_4109));
   NAND3_X1 i_5_4163 (.A1(n_5_1020), .A2(n_5_1019), .A3(n_5_1021), .ZN(n_5_3908));
   INV_X1 i_5_4164 (.A(n_5_3908), .ZN(n_5_3909));
   XNOR2_X1 i_5_4165 (.A(n_5_1591), .B(n_5_1730), .ZN(n_5_3915));
   NAND2_X1 i_5_4166 (.A1(n_5_3915), .A2(n_5_1452), .ZN(n_5_3917));
   NAND3_X1 i_5_1051 (.A1(n_5_3817), .A2(n_5_3818), .A3(n_5_4019), .ZN(n_5_3919));
   NAND3_X1 i_5_1052 (.A1(n_5_3818), .A2(n_5_3817), .A3(n_5_4019), .ZN(n_5_3924));
   INV_X1 i_5_1053 (.A(n_5_3924), .ZN(n_5_3926));
   INV_X1 i_5_4170 (.A(n_5_806), .ZN(n_5_3929));
   NAND3_X1 i_5_4171 (.A1(n_5_436), .A2(n_5_623), .A3(n_5_621), .ZN(n_5_3933));
   NAND2_X1 i_5_4172 (.A1(n_5_623), .A2(n_5_621), .ZN(n_5_3958));
   INV_X1 i_5_4173 (.A(n_5_3958), .ZN(n_5_3962));
   NAND2_X1 i_5_4174 (.A1(n_5_436), .A2(n_5_3962), .ZN(n_5_3980));
   INV_X1 i_5_4175 (.A(n_5_3980), .ZN(n_5_3981));
   NAND2_X1 i_5_2561 (.A1(n_5_4122), .A2(n_5_855), .ZN(n_5_3986));
   NAND2_X1 i_5_4177 (.A1(n_5_917), .A2(n_60), .ZN(n_5_3988));
   INV_X1 i_5_4178 (.A(n_5_855), .ZN(n_5_3992));
   OAI21_X1 i_5_4179 (.A(n_5_3988), .B1(n_5_913), .B2(n_5_3992), .ZN(n_5_4000));
   NAND2_X1 i_5_4180 (.A1(n_5_3664), .A2(n_5_4017), .ZN(n_5_4004));
   NAND2_X1 i_5_4181 (.A1(n_5_3846), .A2(n_5_1006), .ZN(n_5_4014));
   NAND2_X1 i_5_1054 (.A1(n_5_3846), .A2(n_5_1006), .ZN(n_5_4110));
   NAND2_X1 i_5_1084 (.A1(n_5_3664), .A2(n_5_4017), .ZN(n_5_4111));
   INV_X1 i_5_4184 (.A(n_5_4046), .ZN(n_5_4018));
   NAND3_X1 i_5_4185 (.A1(n_5_4109), .A2(n_5_4107), .A3(n_5_4019), .ZN(n_5_4046));
   NAND2_X1 i_5_4186 (.A1(n_5_4019), .A2(n_5_730), .ZN(n_5_4047));
   INV_X1 i_5_4187 (.A(n_5_4047), .ZN(n_5_4112));
   INV_X1 i_5_4188 (.A(n_59), .ZN(n_5_4054));
   NAND2_X1 i_5_4189 (.A1(n_5_724), .A2(n_5_4054), .ZN(n_5_4105));
   INV_X1 i_5_1178 (.A(n_5_4105), .ZN(n_5_4106));
   NAND3_X1 i_5_1185 (.A1(n_5_4517), .A2(n_5_3865), .A3(n_5_4106), .ZN(n_5_4113));
   NAND3_X1 i_5_1097 (.A1(n_5_3775), .A2(n_5_3760), .A3(n_5_3720), .ZN(n_5_4114));
   OR2_X1 i_5_1113 (.A1(n_5_4114), .A2(n_66), .ZN(n_5_4115));
   OR2_X1 i_5_4194 (.A1(n_5_4114), .A2(n_66), .ZN(n_5_4116));
   NAND2_X1 i_5_4195 (.A1(n_5_4114), .A2(n_66), .ZN(n_5_4117));
   NAND2_X1 i_5_4196 (.A1(n_5_4114), .A2(m[5]), .ZN(n_5_4118));
   NAND2_X1 i_5_4197 (.A1(n_5_4114), .A2(m[5]), .ZN(n_5_4119));
   NAND3_X1 i_5_4198 (.A1(n_5_3775), .A2(n_5_3760), .A3(n_5_3720), .ZN(n_5_4120));
   BUF_X1 rt_shieldBuf__2__2__16 (.A(n_5_4187), .Z(n_5_4121));
   INV_X1 i_5_3336 (.A(n_5_913), .ZN(n_5_4122));
   INV_X1 i_5_4200 (.A(n_5_2568), .ZN(n_5_4123));
   NAND2_X1 i_5_4201 (.A1(n_5_570), .A2(n_5_4123), .ZN(n_5_4124));
   INV_X1 i_5_4202 (.A(n_5_4124), .ZN(n_5_4125));
   NAND3_X1 i_5_4203 (.A1(n_5_573), .A2(n_5_3498), .A3(n_5_4125), .ZN(n_5_4126));
   INV_X1 i_5_4204 (.A(n_5_4126), .ZN(n_5_4127));
   INV_X1 i_5_4205 (.A(n_66), .ZN(n_5_4128));
   NAND2_X1 i_5_4206 (.A1(n_5_4699), .A2(n_5_4128), .ZN(n_5_4129));
   INV_X1 i_5_4207 (.A(n_5_4129), .ZN(n_5_4130));
   NAND3_X1 i_5_4208 (.A1(n_5_4697), .A2(n_5_4698), .A3(n_5_4130), .ZN(n_5_4131));
   XNOR2_X1 i_5_4209 (.A(n_5_898), .B(n_5_4000), .ZN(n_5_4132));
   NAND2_X1 i_5_338 (.A1(n_5_4132), .A2(n_5_420), .ZN(n_5_4133));
   NAND3_X1 i_5_3337 (.A1(n_5_1024), .A2(n_5_1025), .A3(n_5_1026), .ZN(n_5_4134));
   NAND2_X1 i_5_3377 (.A1(n_5_4134), .A2(m[8]), .ZN(n_5_4135));
   XNOR2_X1 i_5_4213 (.A(n_5_4134), .B(m[8]), .ZN(n_5_4136));
   OR2_X1 i_5_3384 (.A1(n_5_4134), .A2(m[8]), .ZN(n_5_4137));
   XNOR2_X1 i_5_4215 (.A(n_5_4140), .B(n_60), .ZN(n_5_4138));
   NAND2_X1 i_5_4216 (.A1(n_5_4140), .A2(n_60), .ZN(n_5_4139));
   NAND3_X1 i_5_4217 (.A1(n_5_1024), .A2(n_5_1025), .A3(n_5_1026), .ZN(n_5_4140));
   NAND2_X1 i_5_4220 (.A1(n_5_3933), .A2(n_5_4649), .ZN(n_5_515));
   NAND3_X1 i_5_747 (.A1(n_5_746), .A2(n_5_709), .A3(n_5_911), .ZN(n_5_4141));
   NAND2_X1 i_5_764 (.A1(n_5_786), .A2(n_5_787), .ZN(n_5_4142));
   NAND2_X1 i_5_767 (.A1(n_5_4141), .A2(n_5_4142), .ZN(n_5_4143));
   NAND3_X1 i_5_3385 (.A1(n_5_1016), .A2(n_5_1017), .A3(n_5_1018), .ZN(n_5_4144));
   OR2_X1 i_5_3399 (.A1(n_5_4144), .A2(m[5]), .ZN(n_5_4145));
   NAND2_X1 i_5_3404 (.A1(n_5_4144), .A2(m[5]), .ZN(n_5_4146));
   XNOR2_X1 i_5_4227 (.A(n_5_4144), .B(m[5]), .ZN(n_5_4147));
   NAND2_X1 i_5_4228 (.A1(n_5_4144), .A2(n_66), .ZN(n_5_4148));
   XNOR2_X1 i_5_4229 (.A(n_5_4150), .B(n_66), .ZN(n_5_4149));
   NAND3_X1 i_5_4230 (.A1(n_5_1016), .A2(n_5_1017), .A3(n_5_1018), .ZN(n_5_4150));
   NAND3_X1 i_5_3432 (.A1(n_5_1029), .A2(n_5_3789), .A3(n_5_1030), .ZN(n_5_4151));
   XNOR2_X1 i_5_3433 (.A(n_5_4151), .B(m[10]), .ZN(n_5_4152));
   XNOR2_X1 i_5_3483 (.A(n_5_4151), .B(n_73), .ZN(n_5_4153));
   NAND2_X1 i_5_4234 (.A1(n_5_4151), .A2(n_73), .ZN(n_5_4154));
   NAND3_X1 i_5_4235 (.A1(n_5_1029), .A2(n_5_3789), .A3(n_5_1030), .ZN(n_5_4155));
   NAND2_X1 i_5_4236 (.A1(n_5_3718), .A2(n_5_4119), .ZN(n_5_4156));
   NAND2_X1 i_5_4237 (.A1(n_5_3763), .A2(n_5_3764), .ZN(n_5_4157));
   XNOR2_X1 i_5_4238 (.A(n_5_4156), .B(n_5_4157), .ZN(n_5_4158));
   NAND3_X1 i_5_757 (.A1(n_5_3498), .A2(n_5_573), .A3(n_5_570), .ZN(n_5_4159));
   NAND3_X1 i_5_4240 (.A1(n_5_573), .A2(n_5_3498), .A3(n_5_570), .ZN(n_5_4160));
   NAND2_X1 i_5_4241 (.A1(n_5_4160), .A2(n_5_2568), .ZN(n_5_4161));
   NAND3_X1 i_5_4242 (.A1(n_5_606), .A2(n_5_611), .A3(n_5_605), .ZN(n_5_4162));
   NAND3_X1 i_5_4243 (.A1(n_5_611), .A2(n_5_606), .A3(n_5_605), .ZN(n_5_4163));
   XNOR2_X1 i_5_1128 (.A(n_5_847), .B(n_5_4497), .ZN(n_5_4164));
   NAND2_X1 i_5_1138 (.A1(n_5_4164), .A2(n_5_420), .ZN(n_5_4165));
   NAND3_X1 i_5_4246 (.A1(n_5_4202), .A2(n_5_4393), .A3(n_5_3719), .ZN(n_5_4166));
   INV_X1 i_5_4247 (.A(n_5_4166), .ZN(n_5_4167));
   NAND3_X1 i_5_367 (.A1(n_5_3556), .A2(n_5_4133), .A3(n_5_575), .ZN(n_5_4168));
   XNOR2_X1 i_5_461 (.A(n_5_4168), .B(n_69), .ZN(n_5_4169));
   NAND3_X1 i_5_3544 (.A1(n_5_3556), .A2(n_5_4133), .A3(n_5_575), .ZN(n_5_4170));
   INV_X1 i_5_4251 (.A(n_5_1140), .ZN(n_5_4171));
   INV_X1 i_5_4252 (.A(m[12]), .ZN(n_5_4172));
   XNOR2_X1 i_5_3636 (.A(n_5_3317), .B(n_5_4172), .ZN(n_5_4173));
   XNOR2_X1 i_5_3731 (.A(n_5_1140), .B(n_5_4173), .ZN(n_5_4174));
   NAND2_X1 i_5_4255 (.A1(n_5_732), .A2(n_5_731), .ZN(n_5_4175));
   NAND3_X1 i_5_4256 (.A1(n_5_3505), .A2(n_5_3506), .A3(n_5_3507), .ZN(n_5_4176));
   NAND2_X1 i_5_4257 (.A1(n_5_731), .A2(n_5_732), .ZN(n_5_4177));
   NAND2_X1 i_5_4258 (.A1(n_5_4176), .A2(n_5_4177), .ZN(n_5_4178));
   INV_X1 i_5_4259 (.A(n_5_4178), .ZN(n_5_4179));
   XNOR2_X1 i_5_4260 (.A(n_5_2558), .B(n_5_2363), .ZN(n_5_4180));
   AOI21_X1 i_5_4261 (.A(n_5_2335), .B1(n_5_4180), .B2(n_5_4209), .ZN(n_5_4181));
   NAND2_X1 i_5_4262 (.A1(n_5_923), .A2(n_5_3511), .ZN(n_5_4182));
   NAND2_X1 i_5_4263 (.A1(n_5_3919), .A2(m[4]), .ZN(n_5_4183));
   NAND2_X1 i_5_4264 (.A1(n_5_897), .A2(n_5_420), .ZN(n_5_4184));
   NAND2_X1 i_5_4265 (.A1(n_5_737), .A2(n_5_378), .ZN(n_5_4185));
   NAND2_X1 i_5_4266 (.A1(n_5_3563), .A2(n_5_4649), .ZN(n_5_4186));
   NAND3_X1 i_5_791 (.A1(n_5_4184), .A2(n_5_4185), .A3(n_5_4186), .ZN(n_5_4187));
   NAND3_X1 i_5_773 (.A1(n_5_4424), .A2(n_5_4425), .A3(n_5_4020), .ZN(n_5_4188));
   INV_X1 i_5_4269 (.A(n_5_805), .ZN(n_5_4189));
   NAND2_X1 i_5_4270 (.A1(n_5_804), .A2(n_5_802), .ZN(n_5_4190));
   NAND3_X1 i_5_1166 (.A1(n_5_4189), .A2(n_5_4190), .A3(n_5_3929), .ZN(n_5_4191));
   NAND3_X1 i_5_3576 (.A1(n_5_1019), .A2(n_5_1020), .A3(n_5_1021), .ZN(n_5_4192));
   NAND3_X1 i_5_4273 (.A1(n_5_1020), .A2(n_5_1019), .A3(n_5_1021), .ZN(n_5_4193));
   INV_X1 i_5_4274 (.A(n_5_4193), .ZN(n_5_4194));
   NAND2_X1 i_5_4275 (.A1(n_5_1821), .A2(n_75), .ZN(n_5_4195));
   NAND2_X1 i_5_4276 (.A1(n_5_1705), .A2(n_5_1735), .ZN(n_5_4196));
   NAND3_X1 i_5_4277 (.A1(n_5_1736), .A2(n_5_1754), .A3(n_5_1737), .ZN(n_5_4197));
   NAND2_X1 i_5_4278 (.A1(n_5_1821), .A2(n_75), .ZN(n_5_4198));
   NAND3_X1 i_5_4279 (.A1(n_5_4196), .A2(n_5_4197), .A3(n_5_4198), .ZN(n_5_4199));
   BUF_X1 rt_shieldBuf__2__2__13 (.A(n_50), .Z(n_5_4200));
   XNOR2_X1 i_5_4280 (.A(n_5_2699), .B(n_5_3337), .ZN(n_5_4201));
   NAND2_X1 i_5_1179 (.A1(n_5_4201), .A2(n_5_635), .ZN(n_5_4202));
   NAND2_X1 i_5_465 (.A1(n_5_4165), .A2(n_5_4034), .ZN(n_5_4203));
   XNOR2_X1 i_5_1184 (.A(n_5_4203), .B(n_5_3927), .ZN(n_5_4204));
   OAI22_X1 i_5_4284 (.A1(m[5]), .A2(n_5_4476), .B1(n_5_4203), .B2(m[6]), 
      .ZN(n_5_4205));
   NAND2_X1 i_5_471 (.A1(n_5_4203), .A2(n_5_3185), .ZN(n_5_4206));
   OR2_X1 i_5_472 (.A1(n_5_4203), .A2(n_5_3185), .ZN(n_5_4207));
   NAND2_X1 i_5_3836 (.A1(n_5_4165), .A2(n_5_4034), .ZN(n_5_4208));
   INV_X1 i_5_4288 (.A(n_5_4072), .ZN(n_5_4209));
   XNOR2_X1 i_5_4289 (.A(n_5_4079), .B(n_5_4073), .ZN(n_5_4210));
   INV_X1 i_5_4290 (.A(n_5_4072), .ZN(n_5_4211));
   NAND2_X1 i_5_4291 (.A1(n_5_4210), .A2(n_5_4211), .ZN(n_5_4212));
   NAND3_X1 i_5_525 (.A1(n_5_4348), .A2(n_5_4473), .A3(n_5_3994), .ZN(n_5_4213));
   NAND2_X1 i_5_564 (.A1(n_5_4213), .A2(n_5_4368), .ZN(n_5_4214));
   INV_X1 i_5_583 (.A(n_5_4214), .ZN(n_5_4215));
   NAND2_X1 i_5_4295 (.A1(n_5_4085), .A2(n_5_4065), .ZN(n_5_4216));
   INV_X1 i_5_4296 (.A(n_5_4216), .ZN(n_5_4217));
   OAI21_X1 i_5_4297 (.A(n_5_4217), .B1(n_5_4087), .B2(n_5_4086), .ZN(n_5_4218));
   NAND2_X1 i_5_4298 (.A1(n_5_4078), .A2(n_5_4074), .ZN(n_5_4219));
   INV_X1 i_5_4299 (.A(n_5_4219), .ZN(n_5_4220));
   XNOR2_X1 i_5_4233 (.A(n_5_4356), .B(n_5_3969), .ZN(n_5_4221));
   NAND2_X1 i_5_808 (.A1(n_5_4221), .A2(n_5_188), .ZN(n_5_524));
   XNOR2_X1 i_5_860 (.A(n_5_3886), .B(n_5_3963), .ZN(n_5_4223));
   NAND2_X1 i_5_890 (.A1(n_5_4223), .A2(n_5_188), .ZN(n_5_4663));
   INV_X1 i_5_4304 (.A(m[11]), .ZN(n_5_4224));
   XNOR2_X1 i_5_3851 (.A(n_5_3983), .B(n_5_4224), .ZN(n_5_4225));
   NOR2_X1 i_5_4064 (.A1(n_5_3968), .A2(n_58), .ZN(n_5_4226));
   INV_X1 i_5_4307 (.A(n_5_3968), .ZN(n_5_4227));
   INV_X1 i_5_4308 (.A(n_58), .ZN(n_5_4228));
   NAND2_X1 i_5_4309 (.A1(n_5_4227), .A2(n_5_4228), .ZN(n_5_4229));
   NAND2_X1 i_5_4310 (.A1(n_5_3954), .A2(n_5_4229), .ZN(n_5_4230));
   INV_X1 i_5_4311 (.A(n_5_4230), .ZN(n_5_525));
   NOR2_X1 i_5_4011 (.A1(n_5_4052), .A2(n_65), .ZN(n_5_4232));
   NAND2_X1 i_5_4070 (.A1(n_5_4052), .A2(n_65), .ZN(n_5_4233));
   NAND2_X1 i_5_4314 (.A1(n_5_4052), .A2(n_65), .ZN(n_5_4234));
   INV_X1 i_5_4315 (.A(n_5_4043), .ZN(n_5_4235));
   NOR2_X1 i_5_4316 (.A1(n_5_4052), .A2(n_65), .ZN(n_5_4236));
   OAI21_X1 i_5_4317 (.A(n_5_4234), .B1(n_5_4235), .B2(n_5_4236), .ZN(n_5_4237));
   NAND3_X1 i_5_4318 (.A1(n_5_4107), .A2(n_5_4109), .A3(n_5_4112), .ZN(n_5_4238));
   NAND3_X1 i_5_4319 (.A1(n_5_4109), .A2(n_5_4107), .A3(n_5_4112), .ZN(n_5_4239));
   INV_X1 i_5_4320 (.A(n_5_4239), .ZN(n_5_4240));
   AOI21_X1 i_5_4321 (.A(n_5_4240), .B1(n_5_4182), .B2(n_5_4183), .ZN(n_5_4241));
   XNOR2_X1 i_5_4092 (.A(n_5_3893), .B(n_5_3965), .ZN(n_5_4242));
   NAND2_X1 i_5_4074 (.A1(n_5_4242), .A2(n_5_188), .ZN(n_5_526));
   INV_X1 i_5_4324 (.A(n_65), .ZN(n_5_4243));
   NAND2_X1 i_5_4325 (.A1(n_5_3907), .A2(n_5_4243), .ZN(n_5_4244));
   INV_X1 i_5_4326 (.A(n_5_4244), .ZN(n_5_4245));
   NAND3_X1 i_5_4327 (.A1(n_5_4316), .A2(n_5_4315), .A3(n_5_4245), .ZN(n_5_4246));
   NAND2_X1 i_5_682 (.A1(n_5_4478), .A2(n_5_3869), .ZN(n_5_4248));
   NAND2_X1 i_5_685 (.A1(n_5_3968), .A2(m[4]), .ZN(n_5_4249));
   NAND3_X1 i_5_718 (.A1(n_5_353), .A2(n_5_4248), .A3(n_5_4249), .ZN(n_5_4250));
   NAND2_X1 i_5_4332 (.A1(n_5_4750), .A2(n_5_3877), .ZN(n_5_4251));
   NAND2_X1 i_5_3826 (.A1(n_5_4750), .A2(n_5_3877), .ZN(n_5_4252));
   INV_X1 i_5_524 (.A(n_5_4252), .ZN(n_5_4253));
   NAND2_X1 i_5_3945 (.A1(n_5_4660), .A2(n_60), .ZN(n_5_4254));
   INV_X1 i_5_943 (.A(n_5_4652), .ZN(n_5_4256));
   NAND2_X1 i_5_681 (.A1(n_5_4778), .A2(m[11]), .ZN(n_5_4257));
   XNOR2_X1 i_5_944 (.A(n_5_4778), .B(m[11]), .ZN(n_5_528));
   INV_X1 i_5_3998 (.A(n_5_3863), .ZN(n_5_576));
   XNOR2_X1 i_5_3999 (.A(n_5_4379), .B(n_5_3943), .ZN(n_5_622));
   NAND2_X1 i_5_4343 (.A1(n_5_3968), .A2(m[4]), .ZN(n_5_4262));
   NAND2_X1 i_5_4093 (.A1(n_5_3968), .A2(m[4]), .ZN(n_5_4263));
   INV_X1 i_5_4113 (.A(n_5_4263), .ZN(n_5_4264));
   NAND2_X1 i_5_4346 (.A1(n_5_252), .A2(n_5_226), .ZN(n_5_4265));
   INV_X1 i_5_4347 (.A(n_5_4265), .ZN(n_5_4266));
   NAND2_X1 i_5_836 (.A1(n_5_250), .A2(n_5_4266), .ZN(n_5_531));
   INV_X1 i_5_4350 (.A(n_5_4032), .ZN(n_5_4269));
   NAND2_X1 i_5_983 (.A1(n_5_4024), .A2(n_5_4053), .ZN(n_5_4270));
   NAND2_X1 i_5_1027 (.A1(n_5_4053), .A2(n_5_4024), .ZN(n_5_4271));
   INV_X1 i_5_1028 (.A(n_5_4032), .ZN(n_5_4272));
   INV_X1 i_5_4354 (.A(n_5_4163), .ZN(n_5_4273));
   INV_X1 i_5_4355 (.A(n_5_4021), .ZN(n_5_4274));
   NOR2_X1 i_5_4356 (.A1(n_5_4163), .A2(n_5_4274), .ZN(n_5_4275));
   NAND2_X1 i_5_1082 (.A1(n_5_4791), .A2(n_5_4038), .ZN(n_5_4276));
   NAND3_X1 i_5_1086 (.A1(n_5_4039), .A2(n_5_4035), .A3(n_5_4790), .ZN(n_5_4277));
   NAND2_X1 i_5_1095 (.A1(n_5_4276), .A2(n_5_4277), .ZN(n_5_4278));
   NAND2_X1 i_5_4361 (.A1(n_5_4045), .A2(n_5_4117), .ZN(n_5_4280));
   NAND2_X1 i_5_4362 (.A1(n_5_4049), .A2(n_5_4050), .ZN(n_5_4281));
   NAND3_X1 i_5_4363 (.A1(n_5_4324), .A2(n_5_4280), .A3(n_5_4281), .ZN(n_5_4282));
   OAI21_X1 i_5_1375 (.A(n_5_3941), .B1(n_5_3938), .B2(n_5_3948), .ZN(n_5_4283));
   INV_X1 i_5_4365 (.A(n_5_3964), .ZN(n_5_4284));
   INV_X1 i_5_4366 (.A(n_75), .ZN(n_5_4285));
   NAND2_X1 i_5_4367 (.A1(n_5_4284), .A2(n_5_4285), .ZN(n_5_4286));
   NAND2_X1 i_5_4368 (.A1(n_5_3938), .A2(n_5_3941), .ZN(n_5_4287));
   NAND2_X1 i_5_4369 (.A1(n_5_3948), .A2(n_5_3941), .ZN(n_5_4288));
   NAND3_X1 i_5_3695 (.A1(n_5_4286), .A2(n_5_4287), .A3(n_5_4288), .ZN(n_5_4289));
   INV_X1 i_5_736 (.A(n_5_4246), .ZN(n_5_4290));
   NAND3_X1 i_5_4373 (.A1(n_5_1032), .A2(n_5_4246), .A3(n_5_1373), .ZN(n_5_4292));
   NAND2_X1 i_5_4374 (.A1(n_5_4522), .A2(n_65), .ZN(n_5_4293));
   NAND2_X1 i_5_4375 (.A1(n_5_4292), .A2(n_5_4293), .ZN(n_5_4294));
   NAND2_X1 i_5_821 (.A1(n_5_3888), .A2(n_5_4785), .ZN(n_5_4295));
   NAND2_X1 i_5_1154 (.A1(n_5_4597), .A2(n_5_3880), .ZN(n_5_4296));
   INV_X1 i_5_3972 (.A(n_5_3889), .ZN(n_5_4297));
   NAND3_X1 i_5_4008 (.A1(n_5_4295), .A2(n_5_4296), .A3(n_5_4297), .ZN(n_5_532));
   OR2_X1 i_5_3683 (.A1(n_5_4507), .A2(n_73), .ZN(n_5_4299));
   NAND2_X1 i_5_3752 (.A1(n_5_4507), .A2(n_73), .ZN(n_5_4300));
   XNOR2_X1 i_5_4146 (.A(n_5_4507), .B(n_73), .ZN(n_5_536));
   NOR2_X1 i_5_4383 (.A1(n_5_4461), .A2(m[4]), .ZN(n_5_4302));
   INV_X1 i_5_4384 (.A(n_76), .ZN(n_5_4303));
   XNOR2_X1 i_5_4249 (.A(n_5_3983), .B(n_5_4303), .ZN(n_5_4304));
   XNOR2_X1 i_5_4250 (.A(n_5_4091), .B(n_5_4304), .ZN(n_5_4305));
   NAND3_X1 i_5_1203 (.A1(n_5_4102), .A2(n_5_4088), .A3(n_5_4005), .ZN(n_5_4306));
   XNOR2_X1 i_5_1284 (.A(n_5_4306), .B(n_5_3957), .ZN(n_5_215));
   OR2_X1 i_5_3730 (.A1(n_5_4311), .A2(n_65), .ZN(n_5_4308));
   NAND2_X1 i_5_398 (.A1(n_5_4306), .A2(n_65), .ZN(n_5_4309));
   XNOR2_X1 i_5_3247 (.A(n_5_4306), .B(n_65), .ZN(n_5_216));
   NAND3_X1 i_5_3779 (.A1(n_5_4102), .A2(n_5_4088), .A3(n_5_4005), .ZN(n_5_4311));
   OAI21_X1 i_5_4393 (.A(n_5_4404), .B1(n_5_3883), .B2(n_5_3903), .ZN(n_5_4312));
   NAND2_X1 i_5_4394 (.A1(n_5_429), .A2(n_5_231), .ZN(n_5_4313));
   NAND2_X1 i_5_657 (.A1(n_5_4312), .A2(n_5_4313), .ZN(n_5_4314));
   NAND2_X1 i_5_634 (.A1(n_5_3979), .A2(n_5_197), .ZN(n_5_4315));
   NAND2_X1 i_5_635 (.A1(n_5_3921), .A2(n_5_218), .ZN(n_5_4316));
   NAND2_X1 i_5_3769 (.A1(n_5_3979), .A2(n_5_197), .ZN(n_5_4317));
   INV_X1 i_5_4399 (.A(n_5_3907), .ZN(n_5_4318));
   AOI21_X1 i_5_3793 (.A(n_5_4318), .B1(n_5_3921), .B2(n_5_218), .ZN(n_5_4319));
   NAND2_X1 i_5_3794 (.A1(n_5_4317), .A2(n_5_4319), .ZN(n_5_3873));
   NAND2_X1 i_5_1100 (.A1(n_5_4707), .A2(n_5_4487), .ZN(n_5_4321));
   NAND2_X1 i_5_4114 (.A1(n_5_4044), .A2(n_5_4042), .ZN(n_5_4322));
   AOI21_X1 i_5_4176 (.A(n_5_4045), .B1(n_5_4322), .B2(n_5_4104), .ZN(n_5_4323));
   NAND3_X1 i_5_4405 (.A1(n_5_4325), .A2(n_5_4117), .A3(n_5_4104), .ZN(n_5_4324));
   NAND2_X1 i_5_4406 (.A1(n_5_4044), .A2(n_5_4042), .ZN(n_5_4325));
   NAND3_X1 i_5_4214 (.A1(n_5_3991), .A2(n_5_3990), .A3(n_5_3996), .ZN(n_5_4329));
   NAND2_X1 i_5_4218 (.A1(n_5_616), .A2(n_75), .ZN(n_5_4330));
   XNOR2_X1 i_5_4412 (.A(n_5_3934), .B(n_5_4472), .ZN(n_5_4331));
   NAND2_X1 i_5_935 (.A1(n_5_4331), .A2(n_5_218), .ZN(n_5_4332));
   OAI21_X1 i_5_4414 (.A(n_5_4398), .B1(n_5_4063), .B2(n_5_4064), .ZN(n_5_4333));
   INV_X1 i_5_4415 (.A(n_5_4062), .ZN(n_5_4334));
   OAI21_X1 i_5_4253 (.A(n_5_4398), .B1(n_5_4063), .B2(n_5_4064), .ZN(n_5_4335));
   INV_X1 i_5_4254 (.A(n_5_4062), .ZN(n_5_4336));
   NAND2_X1 i_5_4268 (.A1(n_5_4335), .A2(n_5_4336), .ZN(n_5_4337));
   NAND3_X1 i_5_4282 (.A1(n_5_4730), .A2(n_5_4495), .A3(n_5_3916), .ZN(n_5_4338));
   NAND3_X1 i_5_4136 (.A1(n_5_4730), .A2(n_5_4495), .A3(n_5_3916), .ZN(n_5_4339));
   INV_X1 i_5_4137 (.A(n_5_4339), .ZN(n_5_4340));
   NOR2_X1 i_5_4141 (.A1(n_5_2184), .A2(n_5_4290), .ZN(n_5_4341));
   NAND2_X1 i_5_4167 (.A1(n_5_3967), .A2(n_5_4524), .ZN(n_5_4342));
   NOR2_X1 i_5_4168 (.A1(n_5_4341), .A2(n_5_4342), .ZN(n_5_4343));
   NAND2_X1 i_5_4096 (.A1(n_5_4813), .A2(n_5_218), .ZN(n_5_4346));
   XNOR2_X1 i_5_4292 (.A(n_5_4225), .B(n_5_4057), .ZN(n_5_4347));
   OAI21_X1 i_5_3795 (.A(n_5_4308), .B1(n_5_3987), .B2(n_5_4565), .ZN(n_5_4348));
   AOI21_X1 i_5_4126 (.A(n_5_4559), .B1(n_5_4560), .B2(n_5_4561), .ZN(n_5_219));
   OAI21_X1 i_5_4431 (.A(n_5_3904), .B1(n_5_3905), .B2(n_5_3918), .ZN(n_5_4350));
   NAND2_X1 i_5_4432 (.A1(n_5_4101), .A2(n_59), .ZN(n_5_4351));
   NAND2_X1 i_5_4433 (.A1(n_5_4101), .A2(n_59), .ZN(n_5_4352));
   INV_X1 i_5_4434 (.A(n_5_4352), .ZN(n_5_4353));
   NAND2_X1 i_5_4148 (.A1(n_5_4667), .A2(n_5_3879), .ZN(n_5_539));
   NAND2_X1 i_5_1613 (.A1(n_5_4667), .A2(n_5_3879), .ZN(n_5_4355));
   NAND2_X1 i_5_4285 (.A1(n_5_4435), .A2(n_5_4355), .ZN(n_5_4356));
   NAND3_X1 i_5_4438 (.A1(n_5_4103), .A2(n_5_4013), .A3(n_5_4015), .ZN(n_5_4357));
   NAND2_X1 i_5_4439 (.A1(n_5_4357), .A2(n_61), .ZN(n_5_4358));
   NAND3_X1 i_5_4212 (.A1(n_5_4013), .A2(n_5_4015), .A3(n_5_4103), .ZN(n_5_4359));
   NAND3_X1 i_5_4441 (.A1(n_5_4013), .A2(n_5_4103), .A3(n_5_4015), .ZN(n_5_4360));
   INV_X1 i_5_4442 (.A(n_5_4360), .ZN(n_5_4361));
   NAND2_X1 i_5_4445 (.A1(n_5_4020), .A2(n_5_4036), .ZN(n_5_4364));
   INV_X1 i_5_4446 (.A(n_5_4364), .ZN(n_5_4365));
   NAND3_X1 i_5_4312 (.A1(n_5_4424), .A2(n_5_4425), .A3(n_5_4365), .ZN(n_5_4366));
   OAI21_X1 i_5_4448 (.A(n_5_4131), .B1(n_5_4461), .B2(n_58), .ZN(n_5_4367));
   NAND2_X1 i_5_674 (.A1(n_5_4367), .A2(n_5_4475), .ZN(n_5_4368));
   NAND2_X1 i_5_4182 (.A1(n_5_4258), .A2(n_5_95), .ZN(n_5_546));
   NAND2_X1 i_5_4183 (.A1(n_5_4660), .A2(n_5_3866), .ZN(n_5_578));
   NAND3_X1 i_5_4455 (.A1(n_5_3531), .A2(n_5_185), .A3(n_5_192), .ZN(n_5_4373));
   INV_X1 i_5_4456 (.A(n_5_4373), .ZN(n_5_4374));
   INV_X1 i_5_4457 (.A(n_5_3953), .ZN(n_5_4375));
   NAND2_X1 i_5_4458 (.A1(n_5_4374), .A2(n_5_4375), .ZN(n_5_4376));
   INV_X1 i_5_4459 (.A(n_5_3952), .ZN(n_5_4377));
   NAND2_X1 i_5_4460 (.A1(n_5_4373), .A2(n_5_4377), .ZN(n_5_4378));
   NAND2_X1 i_5_4340 (.A1(n_5_4376), .A2(n_5_4378), .ZN(n_5_4379));
   NAND2_X1 i_5_4219 (.A1(n_5_4329), .A2(n_5_4330), .ZN(n_5_579));
   NAND2_X1 i_5_4224 (.A1(n_5_3989), .A2(n_5_4358), .ZN(n_5_581));
   INV_X1 i_5_4465 (.A(n_5_4100), .ZN(n_5_4383));
   NAND2_X1 i_5_4466 (.A1(n_5_4094), .A2(n_5_4096), .ZN(n_5_4384));
   NAND2_X1 i_5_4467 (.A1(n_5_4383), .A2(n_5_4384), .ZN(n_5_4385));
   NAND2_X1 i_5_4468 (.A1(n_5_4025), .A2(n_5_4029), .ZN(n_5_4386));
   INV_X1 i_5_4469 (.A(n_5_4386), .ZN(n_5_4387));
   NAND2_X1 i_5_4470 (.A1(n_5_4026), .A2(n_5_4387), .ZN(n_5_4388));
   INV_X1 i_5_4471 (.A(n_5_4388), .ZN(n_5_4389));
   XNOR2_X1 i_5_4474 (.A(n_5_4089), .B(n_5_4097), .ZN(n_5_4392));
   NAND2_X1 i_5_4192 (.A1(n_5_4392), .A2(n_5_4017), .ZN(n_5_4393));
   NAND3_X1 i_5_4476 (.A1(n_5_4082), .A2(n_5_4083), .A3(n_5_4084), .ZN(n_5_4394));
   INV_X1 i_5_4477 (.A(n_69), .ZN(n_5_4395));
   NAND2_X1 i_5_4478 (.A1(n_5_4084), .A2(n_5_4395), .ZN(n_5_4396));
   INV_X1 i_5_4479 (.A(n_5_4396), .ZN(n_5_4397));
   NAND3_X1 i_5_4302 (.A1(n_5_4082), .A2(n_5_4083), .A3(n_5_4397), .ZN(n_5_4398));
   NAND3_X1 i_5_4481 (.A1(n_5_4107), .A2(n_5_4109), .A3(n_5_4019), .ZN(n_5_4399));
   NAND2_X1 i_5_4193 (.A1(n_5_4399), .A2(n_58), .ZN(n_5_4400));
   NAND2_X1 i_5_4210 (.A1(n_5_4715), .A2(n_66), .ZN(n_5_4401));
   XNOR2_X1 i_5_4244 (.A(n_5_4715), .B(n_5_3898), .ZN(n_5_4402));
   XNOR2_X1 i_5_4485 (.A(n_5_4715), .B(n_5_3940), .ZN(n_5_4403));
   NAND2_X1 i_5_4486 (.A1(n_5_4715), .A2(m[5]), .ZN(n_5_4404));
   NAND3_X1 i_5_4377 (.A1(n_5_4011), .A2(n_5_4012), .A3(n_5_4010), .ZN(n_5_616));
   NAND3_X1 i_5_4488 (.A1(n_5_4011), .A2(n_5_4012), .A3(n_5_4010), .ZN(n_5_4406));
   INV_X1 i_5_4489 (.A(n_5_4406), .ZN(n_5_4407));
   NAND2_X1 i_5_4490 (.A1(n_5_4522), .A2(n_5_3866), .ZN(n_5_4408));
   NAND2_X1 i_5_4493 (.A1(n_5_4522), .A2(n_5_3866), .ZN(n_5_625));
   NAND3_X1 i_5_697 (.A1(n_5_518), .A2(n_5_3928), .A3(n_5_459), .ZN(n_5_4412));
   NAND3_X1 i_5_717 (.A1(n_5_4586), .A2(n_5_4412), .A3(n_5_218), .ZN(n_5_4413));
   NAND2_X1 i_5_4221 (.A1(m[9]), .A2(n_5_4686), .ZN(n_5_4414));
   NAND2_X1 i_5_1187 (.A1(n_5_4271), .A2(n_5_4272), .ZN(n_5_4415));
   NAND2_X1 i_5_4335 (.A1(n_5_4023), .A2(n_5_4270), .ZN(n_5_4416));
   AOI22_X1 i_5_4337 (.A1(n_5_4271), .A2(n_5_4272), .B1(n_5_4686), .B2(m[9]), 
      .ZN(n_5_4417));
   NAND2_X1 i_5_4338 (.A1(n_5_4416), .A2(n_5_4417), .ZN(n_5_626));
   XNOR2_X1 i_5_4245 (.A(n_5_3882), .B(n_5_4402), .ZN(n_5_646));
   NAND3_X1 i_5_4305 (.A1(n_5_878), .A2(n_5_3959), .A3(n_5_196), .ZN(n_5_4422));
   NAND2_X1 i_5_4323 (.A1(n_5_4422), .A2(n_73), .ZN(n_5_4423));
   NAND2_X1 i_5_4341 (.A1(n_5_4305), .A2(n_5_4017), .ZN(n_5_4424));
   NAND2_X1 i_5_4351 (.A1(n_5_4347), .A2(n_5_1006), .ZN(n_5_4425));
   NAND2_X1 i_5_3347 (.A1(n_5_4305), .A2(n_5_4017), .ZN(n_5_4426));
   NAND2_X1 i_5_3380 (.A1(n_5_4347), .A2(n_5_1006), .ZN(n_5_4427));
   NAND3_X1 i_5_3487 (.A1(n_5_4426), .A2(n_5_4427), .A3(n_5_4020), .ZN(n_5_4428));
   NAND2_X1 i_5_4514 (.A1(n_5_159), .A2(n_5_160), .ZN(n_5_4429));
   OAI21_X1 i_5_4515 (.A(n_5_4779), .B1(n_5_4781), .B2(n_5_4780), .ZN(n_5_4430));
   NAND2_X1 i_5_4516 (.A1(n_5_4429), .A2(n_5_4430), .ZN(n_5_4431));
   NAND2_X1 i_5_3995 (.A1(n_5_4665), .A2(m[10]), .ZN(n_5_4432));
   NAND2_X1 i_5_4301 (.A1(n_5_4251), .A2(n_5_3887), .ZN(n_5_4433));
   NAND2_X1 i_5_4408 (.A1(n_5_4748), .A2(m[9]), .ZN(n_5_4434));
   NAND3_X1 i_5_4436 (.A1(n_5_4432), .A2(n_5_4433), .A3(n_5_4434), .ZN(n_5_4435));
   NAND3_X1 i_5_646 (.A1(n_5_3972), .A2(n_5_3973), .A3(n_5_3906), .ZN(n_5_4436));
   NAND3_X1 i_5_4423 (.A1(n_5_3971), .A2(n_5_4520), .A3(n_5_3950), .ZN(n_5_4437));
   NAND3_X1 i_5_4424 (.A1(n_5_3972), .A2(n_5_3973), .A3(n_5_3906), .ZN(n_5_4438));
   NAND2_X1 i_5_4512 (.A1(n_5_4437), .A2(n_5_4438), .ZN(n_5_647));
   NAND3_X1 i_5_4525 (.A1(n_5_4077), .A2(n_5_4075), .A3(n_5_4076), .ZN(n_5_4440));
   NAND2_X1 i_5_4526 (.A1(n_48), .A2(n_60), .ZN(n_5_4441));
   NAND3_X1 i_5_4527 (.A1(n_5_4075), .A2(n_5_4076), .A3(n_5_4077), .ZN(n_5_4442));
   NAND2_X1 i_5_4528 (.A1(n_48), .A2(n_60), .ZN(n_5_4443));
   NAND2_X1 i_5_4529 (.A1(n_5_4442), .A2(n_5_4443), .ZN(n_5_4444));
   NAND2_X1 i_5_4530 (.A1(n_5_4033), .A2(n_5_4027), .ZN(n_5_4445));
   NAND2_X1 i_5_4531 (.A1(n_5_4028), .A2(n_5_4241), .ZN(n_5_4446));
   NAND2_X1 i_5_4532 (.A1(n_5_4445), .A2(n_5_4446), .ZN(n_5_876));
   INV_X1 i_5_4533 (.A(n_5_4449), .ZN(n_5_4448));
   NAND3_X1 i_5_4169 (.A1(n_5_4346), .A2(n_5_4806), .A3(n_5_3906), .ZN(n_5_4449));
   NAND2_X1 i_5_4535 (.A1(n_5_3906), .A2(n_5_3868), .ZN(n_5_4450));
   INV_X1 i_5_4536 (.A(n_5_4450), .ZN(n_5_4451));
   NAND3_X1 i_5_4537 (.A1(n_5_4806), .A2(n_5_4346), .A3(n_5_4451), .ZN(n_5_4452));
   NAND2_X1 i_5_4232 (.A1(n_5_4022), .A2(n_5_4031), .ZN(n_5_4453));
   INV_X1 i_5_4300 (.A(n_5_4453), .ZN(n_5_4454));
   NAND2_X1 i_5_4540 (.A1(n_5_4066), .A2(n_5_4080), .ZN(n_5_4455));
   NAND3_X1 i_5_4541 (.A1(n_5_4066), .A2(n_5_4080), .A3(n_5_4081), .ZN(n_5_4456));
   NAND3_X1 i_5_4542 (.A1(n_5_4007), .A2(n_5_4056), .A3(n_5_4006), .ZN(n_5_4457));
   XNOR2_X1 i_5_4095 (.A(n_5_4457), .B(n_58), .ZN(n_5_4458));
   NAND2_X1 i_5_4544 (.A1(n_5_4457), .A2(m[4]), .ZN(n_5_256));
   XNOR2_X1 i_5_4545 (.A(n_5_4457), .B(m[4]), .ZN(n_5_4460));
   NAND3_X1 i_5_4546 (.A1(n_5_4007), .A2(n_5_4056), .A3(n_5_4006), .ZN(n_5_4461));
   NAND3_X1 i_5_4548 (.A1(n_5_4463), .A2(n_5_4464), .A3(n_5_4067), .ZN(n_5_4462));
   NAND2_X1 i_5_4549 (.A1(n_5_4070), .A2(n_5_4069), .ZN(n_5_4463));
   NAND2_X1 i_5_4550 (.A1(n_5_4071), .A2(n_5_4068), .ZN(n_5_4464));
   NAND2_X1 i_5_4551 (.A1(n_5_4070), .A2(n_5_4069), .ZN(n_5_4465));
   INV_X1 i_5_4552 (.A(n_5_4068), .ZN(n_5_4466));
   NAND2_X1 i_5_4553 (.A1(n_5_4067), .A2(n_5_4466), .ZN(n_5_4467));
   INV_X1 i_5_4554 (.A(n_5_4067), .ZN(n_5_4468));
   OAI21_X1 i_5_4555 (.A(n_5_4467), .B1(n_5_4071), .B2(n_5_4468), .ZN(n_5_4469));
   NAND2_X1 i_5_4556 (.A1(n_5_4465), .A2(n_5_4469), .ZN(n_5_4470));
   INV_X1 i_5_4557 (.A(n_5_4470), .ZN(n_5_4471));
   XNOR2_X1 i_5_4558 (.A(n_5_4703), .B(m[5]), .ZN(n_5_4472));
   NAND2_X1 i_5_4559 (.A1(n_5_4703), .A2(n_66), .ZN(n_5_4473));
   XNOR2_X1 i_5_4286 (.A(n_5_4703), .B(n_66), .ZN(n_5_4474));
   NAND2_X1 i_5_4561 (.A1(n_5_4703), .A2(n_66), .ZN(n_5_4475));
   NAND3_X1 i_5_4271 (.A1(n_5_4697), .A2(n_5_4698), .A3(n_5_4699), .ZN(n_5_4476));
   NAND2_X1 i_5_4563 (.A1(n_5_3881), .A2(n_5_4452), .ZN(n_5_4477));
   INV_X1 i_5_4564 (.A(n_5_4477), .ZN(n_5_4478));
   XNOR2_X1 i_5_4380 (.A(n_5_3998), .B(n_5_4474), .ZN(n_5_4479));
   NAND2_X1 i_5_4413 (.A1(n_5_4479), .A2(n_5_197), .ZN(n_5_4480));
   NAND2_X1 i_5_4567 (.A1(n_5_4108), .A2(n_55), .ZN(n_5_4481));
   OAI21_X1 i_5_4568 (.A(n_5_4095), .B1(n_5_4108), .B2(n_55), .ZN(n_5_4482));
   NAND2_X1 i_5_4569 (.A1(n_5_4108), .A2(n_55), .ZN(n_5_4483));
   NOR2_X1 i_5_4570 (.A1(n_5_4090), .A2(n_5_4098), .ZN(n_5_4484));
   NAND3_X1 i_5_4117 (.A1(n_5_4775), .A2(n_5_4774), .A3(n_5_515), .ZN(n_5_4486));
   NAND2_X1 i_5_4139 (.A1(n_5_4486), .A2(n_76), .ZN(n_5_4487));
   INV_X1 i_5_4574 (.A(n_5_90), .ZN(n_5_4488));
   XNOR2_X1 i_5_4575 (.A(n_5_94), .B(n_5_4488), .ZN(n_5_4489));
   INV_X1 i_5_4576 (.A(n_5_3855), .ZN(n_5_4490));
   OAI22_X1 i_5_4577 (.A1(n_5_4489), .A2(n_5_4490), .B1(n_5_3855), .B2(n_5_90), 
      .ZN(n_5_4670));
   NAND2_X1 i_5_116 (.A1(n_5_4523), .A2(m[8]), .ZN(n_5_4492));
   NAND2_X1 i_5_726 (.A1(n_5_4594), .A2(n_5_4492), .ZN(n_5_4493));
   NAND2_X1 i_5_4487 (.A1(n_5_3681), .A2(n_5_197), .ZN(n_5_4495));
   NAND3_X1 i_5_4281 (.A1(n_5_4110), .A2(n_5_4111), .A3(n_5_4016), .ZN(n_5_4496));
   XNOR2_X1 i_5_4283 (.A(n_5_4496), .B(n_5_4048), .ZN(n_5_4497));
   INV_X1 i_5_4585 (.A(n_5_4499), .ZN(n_5_4498));
   NAND3_X1 i_5_4586 (.A1(n_5_4110), .A2(n_5_4111), .A3(n_5_4016), .ZN(n_5_4499));
   NAND3_X1 i_5_742 (.A1(n_5_3920), .A2(n_5_4413), .A3(n_5_3910), .ZN(n_5_4500));
   NAND3_X1 i_5_775 (.A1(n_5_3920), .A2(n_5_4413), .A3(n_5_3910), .ZN(n_5_4501));
   INV_X1 i_5_1182 (.A(n_5_4500), .ZN(n_5_294));
   AND2_X1 i_5_3630 (.A1(n_5_4501), .A2(n_5_3185), .ZN(n_5_4503));
   XNOR2_X1 i_5_4010 (.A(n_5_4500), .B(n_5_3949), .ZN(n_5_4504));
   NAND2_X1 i_5_4592 (.A1(n_5_3736), .A2(n_5_4041), .ZN(n_5_4505));
   INV_X1 i_5_4593 (.A(n_5_3808), .ZN(n_5_4506));
   NAND3_X1 i_5_3637 (.A1(n_5_4001), .A2(n_5_4002), .A3(n_5_4003), .ZN(n_5_4507));
   NAND3_X1 i_5_3672 (.A1(n_5_4001), .A2(n_5_4002), .A3(n_5_4003), .ZN(n_5_4508));
   INV_X1 i_5_3873 (.A(n_5_4508), .ZN(n_5_649));
   INV_X1 i_5_4597 (.A(n_5_4099), .ZN(n_5_4510));
   NAND2_X1 i_5_4598 (.A1(n_5_4092), .A2(n_5_4093), .ZN(n_5_4511));
   XNOR2_X1 i_5_4599 (.A(n_5_4511), .B(n_5_4099), .ZN(n_5_4512));
   AOI21_X1 i_5_3996 (.A(n_5_4256), .B1(n_5_3944), .B2(n_5_3942), .ZN(n_5_4513));
   AOI21_X1 i_5_3997 (.A(n_5_3939), .B1(n_5_3951), .B2(n_5_4513), .ZN(n_5_4514));
   AOI21_X1 i_5_4443 (.A(n_5_4256), .B1(n_5_3944), .B2(n_5_3942), .ZN(n_5_4515));
   XNOR2_X1 i_5_4329 (.A(n_5_4051), .B(n_5_4030), .ZN(n_5_4516));
   NAND2_X1 i_5_4330 (.A1(n_5_4516), .A2(n_5_378), .ZN(n_5_4517));
   OAI21_X1 i_5_4605 (.A(n_5_3904), .B1(n_5_3905), .B2(n_5_3918), .ZN(n_5_4518));
   OAI21_X1 i_5_4344 (.A(n_5_3904), .B1(n_5_3905), .B2(n_5_3918), .ZN(n_5_4519));
   NAND2_X1 i_5_4348 (.A1(n_5_4519), .A2(m[0]), .ZN(n_5_4520));
   NAND3_X1 i_5_721 (.A1(n_5_4315), .A2(n_5_4316), .A3(n_5_3907), .ZN(n_5_291));
   NAND3_X1 i_5_4609 (.A1(n_5_4315), .A2(n_5_4316), .A3(n_5_3907), .ZN(n_5_4522));
   INV_X1 i_5_740 (.A(n_5_291), .ZN(n_5_316));
   NAND2_X1 i_5_4611 (.A1(n_5_4522), .A2(n_65), .ZN(n_5_4524));
   INV_X1 i_5_4239 (.A(n_5_3970), .ZN(n_5_4526));
   NAND2_X1 i_5_4267 (.A1(n_5_4350), .A2(m[0]), .ZN(n_5_4527));
   NAND2_X1 i_5_4615 (.A1(n_5_4350), .A2(m[0]), .ZN(n_5_4528));
   INV_X1 i_5_4616 (.A(n_5_4528), .ZN(n_5_4529));
   INV_X1 i_5_4617 (.A(n_5_3867), .ZN(n_5_4530));
   OAI21_X1 i_5_4618 (.A(n_5_4529), .B1(n_5_3970), .B2(n_5_4530), .ZN(n_5_4531));
   NAND3_X1 i_5_4000 (.A1(n_5_4059), .A2(n_5_4060), .A3(n_5_4061), .ZN(n_5_678));
   NAND3_X1 i_5_4620 (.A1(n_5_4059), .A2(n_5_4060), .A3(n_5_4061), .ZN(n_5_4533));
   INV_X1 i_5_4621 (.A(n_5_4533), .ZN(n_5_4534));
   NAND2_X1 i_5_4045 (.A1(n_5_4372), .A2(n_5_3975), .ZN(n_5_4538));
   INV_X1 i_5_4055 (.A(n_5_4538), .ZN(n_5_4671));
   INV_X1 i_5_4628 (.A(n_5_4547), .ZN(n_5_684));
   NAND2_X1 i_5_4629 (.A1(n_5_157), .A2(n_5_158), .ZN(n_5_692));
   NAND3_X1 i_5_4589 (.A1(n_5_163), .A2(n_5_162), .A3(n_5_181), .ZN(n_5_3890));
   NAND2_X1 i_5_4637 (.A1(n_5_4668), .A2(n_5_4691), .ZN(n_5_4548));
   NAND2_X1 i_5_4638 (.A1(m[11]), .A2(n_5_293), .ZN(n_5_4549));
   NAND2_X1 i_5_4364 (.A1(n_5_279), .A2(n_5_188), .ZN(n_5_4553));
   NAND2_X1 i_5_4370 (.A1(n_5_568), .A2(n_5_95), .ZN(n_5_4554));
   NAND3_X1 i_5_4381 (.A1(n_5_4553), .A2(n_5_4554), .A3(n_5_227), .ZN(n_5_4672));
   INV_X1 i_5_4649 (.A(n_5_4113), .ZN(n_5_4559));
   NAND2_X1 i_5_4650 (.A1(n_5_620), .A2(n_5_723), .ZN(n_5_4560));
   NAND2_X1 i_5_4651 (.A1(n_5_4566), .A2(n_59), .ZN(n_5_4561));
   INV_X1 i_5_4190 (.A(n_5_4113), .ZN(n_5_4562));
   NAND2_X1 i_5_4191 (.A1(n_5_723), .A2(n_5_620), .ZN(n_5_4563));
   NAND2_X1 i_5_4211 (.A1(n_5_4566), .A2(n_59), .ZN(n_5_4564));
   AOI21_X1 i_5_4225 (.A(n_5_4562), .B1(n_5_4563), .B2(n_5_4564), .ZN(n_5_4565));
   NAND3_X1 i_5_4371 (.A1(n_5_4517), .A2(n_5_3865), .A3(n_5_724), .ZN(n_5_4566));
   NAND2_X1 i_5_4387 (.A1(n_5_503), .A2(n_5_522), .ZN(n_5_432));
   INV_X1 i_5_4658 (.A(m[2]), .ZN(n_5_4568));
   NAND2_X1 i_5_4659 (.A1(n_5_724), .A2(n_5_4568), .ZN(n_5_4569));
   INV_X1 i_5_4660 (.A(n_5_4569), .ZN(n_5_4570));
   NAND3_X1 i_5_4388 (.A1(n_5_3865), .A2(n_5_4517), .A3(n_5_4570), .ZN(n_5_443));
   OAI21_X1 i_5_3634 (.A(n_5_4483), .B1(n_5_4482), .B2(n_5_4484), .ZN(n_5_4573));
   NAND2_X1 i_5_4664 (.A1(n_5_4506), .A2(n_5_4505), .ZN(n_5_4574));
   NAND3_X1 i_5_4665 (.A1(n_5_3808), .A2(n_5_3736), .A3(n_5_3682), .ZN(n_5_4575));
   NAND2_X1 i_5_4499 (.A1(n_5_4574), .A2(n_5_4575), .ZN(n_5_700));
   NAND2_X1 i_5_4667 (.A1(n_5_4660), .A2(m[8]), .ZN(n_5_4577));
   INV_X1 i_5_550 (.A(n_5_4651), .ZN(n_5_4673));
   INV_X1 i_5_4670 (.A(n_5_4580), .ZN(n_5_429));
   NAND3_X1 i_5_4671 (.A1(n_5_4712), .A2(n_5_4711), .A3(n_5_4627), .ZN(n_5_4580));
   NAND2_X1 i_5_4672 (.A1(n_5_4627), .A2(n_5_231), .ZN(n_5_4581));
   INV_X1 i_5_4673 (.A(n_5_4581), .ZN(n_5_4582));
   NAND3_X1 i_5_4674 (.A1(n_5_4712), .A2(n_5_4711), .A3(n_5_4582), .ZN(n_5_4583));
   NAND2_X1 i_5_4024 (.A1(n_5_518), .A2(n_5_459), .ZN(n_5_4584));
   INV_X1 i_5_4026 (.A(n_5_475), .ZN(n_5_4585));
   NAND2_X1 i_5_4038 (.A1(n_5_4584), .A2(n_5_4585), .ZN(n_5_4586));
   XNOR2_X1 i_5_3667 (.A(n_5_3864), .B(n_5_4152), .ZN(n_5_4587));
   NAND2_X1 i_5_3719 (.A1(n_5_4587), .A2(n_5_1006), .ZN(n_5_4588));
   NAND3_X1 i_5_4062 (.A1(n_5_4620), .A2(n_5_4621), .A3(n_5_4622), .ZN(n_5_4674));
   OR2_X1 i_5_222 (.A1(n_5_4674), .A2(n_66), .ZN(n_5_4675));
   NAND2_X1 i_5_484 (.A1(n_5_4679), .A2(n_66), .ZN(n_5_4676));
   NAND2_X1 i_5_4199 (.A1(n_5_4674), .A2(m[5]), .ZN(n_5_4677));
   OR2_X1 i_5_4231 (.A1(n_5_4674), .A2(m[5]), .ZN(n_5_4678));
   NAND3_X1 i_5_4287 (.A1(n_5_4620), .A2(n_5_4621), .A3(n_5_4622), .ZN(n_5_4679));
   NAND2_X1 i_5_4686 (.A1(n_5_4636), .A2(n_5_4637), .ZN(n_5_4680));
   NAND2_X1 i_5_4687 (.A1(n_5_4642), .A2(n_5_197), .ZN(n_5_4681));
   NAND3_X1 i_5_4306 (.A1(n_5_4680), .A2(n_5_4681), .A3(n_5_4627), .ZN(n_5_4682));
   XNOR2_X1 i_5_4689 (.A(n_5_4644), .B(n_5_381), .ZN(n_5_4683));
   INV_X1 i_5_4690 (.A(n_5_4644), .ZN(n_5_4684));
   XNOR2_X1 i_5_4691 (.A(n_5_381), .B(n_5_4684), .ZN(n_5_4685));
   NAND2_X1 i_5_4447 (.A1(n_5_4656), .A2(n_5_4657), .ZN(n_5_4686));
   NAND2_X1 i_5_4693 (.A1(n_5_4657), .A2(n_5_4656), .ZN(n_5_4687));
   NAND2_X1 i_5_4694 (.A1(n_5_4687), .A2(m[9]), .ZN(n_5_4688));
   NAND2_X1 i_5_4631 (.A1(n_5_4261), .A2(n_5_197), .ZN(n_5_4689));
   NAND2_X1 i_5_4632 (.A1(n_5_4631), .A2(n_5_218), .ZN(n_5_4690));
   NAND2_X1 i_5_4452 (.A1(n_5_4631), .A2(n_5_218), .ZN(n_5_701));
   NAND3_X1 i_5_4389 (.A1(n_5_4659), .A2(n_5_4658), .A3(n_5_4653), .ZN(n_5_4694));
   NAND3_X1 i_5_4701 (.A1(n_5_4659), .A2(n_5_4658), .A3(n_5_4653), .ZN(n_5_4695));
   INV_X1 i_5_4702 (.A(n_5_4695), .ZN(n_5_4696));
   NAND2_X1 i_5_4398 (.A1(n_5_4222), .A2(n_5_378), .ZN(n_5_4697));
   NAND2_X1 i_5_4403 (.A1(n_5_4655), .A2(n_5_420), .ZN(n_5_4698));
   NAND2_X1 i_5_4705 (.A1(n_5_4694), .A2(n_5_4649), .ZN(n_5_4699));
   NAND2_X1 i_5_4517 (.A1(n_5_4655), .A2(n_5_420), .ZN(n_5_4700));
   NAND2_X1 i_5_4708 (.A1(n_5_4694), .A2(n_5_4649), .ZN(n_5_4702));
   NAND3_X1 i_5_4560 (.A1(n_5_4700), .A2(n_5_4600), .A3(n_5_4702), .ZN(n_5_4703));
   INV_X1 i_5_4710 (.A(n_5_4589), .ZN(n_5_4704));
   NAND3_X1 i_5_4711 (.A1(n_5_4775), .A2(n_5_4774), .A3(n_5_515), .ZN(n_5_4589));
   NAND2_X1 i_5_4712 (.A1(n_5_515), .A2(n_5_4645), .ZN(n_5_4705));
   INV_X1 i_5_4334 (.A(n_5_4705), .ZN(n_5_4706));
   NAND3_X1 i_5_4352 (.A1(n_5_4775), .A2(n_5_4774), .A3(n_5_4706), .ZN(n_5_4707));
   NAND2_X1 i_5_4416 (.A1(n_5_4673), .A2(n_5_4626), .ZN(n_5_4709));
   NAND2_X1 i_5_4421 (.A1(n_5_1031), .A2(n_5_4709), .ZN(n_5_465));
   NAND2_X1 i_5_4718 (.A1(n_5_4636), .A2(n_5_4637), .ZN(n_5_4711));
   NAND2_X1 i_5_4719 (.A1(n_5_4642), .A2(n_5_197), .ZN(n_5_4712));
   NAND2_X1 i_5_4404 (.A1(n_5_4636), .A2(n_5_4637), .ZN(n_5_4713));
   NAND2_X1 i_5_4410 (.A1(n_5_4642), .A2(n_5_197), .ZN(n_5_4714));
   NAND3_X1 i_5_4484 (.A1(n_5_4713), .A2(n_5_4714), .A3(n_5_4627), .ZN(n_5_4715));
   NAND3_X1 i_5_4496 (.A1(n_5_347), .A2(n_5_526), .A3(n_5_132), .ZN(n_5_702));
   XNOR2_X1 i_5_4085 (.A(n_5_702), .B(n_5_3185), .ZN(n_5_4718));
   NAND3_X1 i_5_4418 (.A1(n_5_347), .A2(n_5_526), .A3(n_5_132), .ZN(n_5_711));
   AOI21_X1 i_5_4480 (.A(n_5_4646), .B1(n_5_4648), .B2(n_5_4647), .ZN(n_5_716));
   NAND2_X1 i_5_4353 (.A1(n_5_4648), .A2(n_5_4647), .ZN(n_5_728));
   INV_X1 i_5_4357 (.A(n_5_4646), .ZN(n_5_739));
   XNOR2_X1 i_5_4336 (.A(n_5_4671), .B(n_5_4809), .ZN(n_5_3705));
   NAND2_X1 i_5_4138 (.A1(n_5_4634), .A2(n_5_4633), .ZN(n_5_4728));
   NAND2_X1 i_5_4322 (.A1(n_5_4633), .A2(n_5_4632), .ZN(n_5_4729));
   NAND3_X1 i_5_4328 (.A1(n_5_4728), .A2(n_5_4729), .A3(n_5_218), .ZN(n_5_4730));
   NAND3_X1 i_5_4088 (.A1(n_5_4663), .A2(n_5_4639), .A3(n_5_4640), .ZN(n_5_4731));
   XNOR2_X1 i_5_660 (.A(n_5_4731), .B(m[9]), .ZN(n_5_4732));
   NOR2_X1 i_5_4115 (.A1(n_5_4731), .A2(n_55), .ZN(n_5_3706));
   XNOR2_X1 i_5_4407 (.A(n_5_4731), .B(n_55), .ZN(n_5_4734));
   NAND3_X1 i_5_4116 (.A1(n_5_4663), .A2(n_5_4639), .A3(n_5_4640), .ZN(n_5_3856));
   NAND2_X1 i_5_3767 (.A1(n_5_159), .A2(n_5_160), .ZN(n_5_749));
   NAND2_X1 i_5_4461 (.A1(n_5_159), .A2(n_5_160), .ZN(n_5_821));
   NAND2_X1 i_5_4472 (.A1(n_5_3874), .A2(n_5_821), .ZN(n_5_1031));
   NAND3_X1 i_5_4716 (.A1(n_5_647), .A2(n_5_355), .A3(n_5_333), .ZN(n_5_1032));
   NAND2_X1 i_5_4717 (.A1(n_5_327), .A2(n_5_354), .ZN(n_5_1373));
   NAND3_X1 i_5_4607 (.A1(n_5_647), .A2(n_5_333), .A3(n_5_355), .ZN(n_5_1374));
   NAND2_X1 i_5_4723 (.A1(n_5_327), .A2(n_5_354), .ZN(n_5_1382));
   NAND2_X1 i_5_4734 (.A1(n_5_1374), .A2(n_5_1382), .ZN(n_5_2184));
   XNOR2_X1 i_5_4494 (.A(n_5_536), .B(n_5_4371), .ZN(n_5_3353));
   NAND2_X1 i_5_4579 (.A1(n_5_3353), .A2(n_5_197), .ZN(n_5_3531));
   INV_X1 i_5_4379 (.A(n_75), .ZN(n_5_3632));
   XNOR2_X1 i_5_4727 (.A(n_5_616), .B(n_5_3632), .ZN(n_5_3639));
   XNOR2_X1 i_5_4728 (.A(n_5_3639), .B(n_5_372), .ZN(n_5_3681));
   INV_X1 i_5_4735 (.A(m[11]), .ZN(n_5_3707));
   NAND2_X1 i_5_4736 (.A1(n_5_515), .A2(n_5_3707), .ZN(n_5_3708));
   INV_X1 i_5_4739 (.A(n_5_3708), .ZN(n_5_3709));
   NAND3_X1 i_5_4740 (.A1(n_5_4774), .A2(n_5_4775), .A3(n_5_3709), .ZN(n_5_3710));
   NAND2_X1 i_5_4741 (.A1(n_5_649), .A2(n_5_251), .ZN(n_5_3806));
   NAND2_X1 i_5_4345 (.A1(n_5_3710), .A2(n_5_3806), .ZN(n_5_3807));
   INV_X1 i_5_4729 (.A(n_5_684), .ZN(n_5_3809));
   INV_X1 i_5_4743 (.A(n_5_692), .ZN(n_5_3871));
   AOI21_X1 i_5_4744 (.A(n_5_4763), .B1(n_5_4764), .B2(n_5_4765), .ZN(n_5_3872));
   OAI21_X1 i_5_4547 (.A(n_5_3809), .B1(n_5_3871), .B2(n_5_3872), .ZN(n_5_3874));
   NAND2_X1 i_5_4142 (.A1(n_5_486), .A2(n_5_476), .ZN(n_5_3875));
   XNOR2_X1 i_5_4223 (.A(n_5_497), .B(n_5_678), .ZN(n_5_3876));
   OAI21_X1 i_5_4248 (.A(n_5_3875), .B1(n_5_3876), .B2(n_5_486), .ZN(n_5_3878));
   NAND3_X1 i_5_4422 (.A1(n_5_4625), .A2(n_5_4628), .A3(n_5_183), .ZN(n_5_3930));
   INV_X1 i_5_4738 (.A(n_69), .ZN(n_5_3895));
   NAND2_X1 i_5_4746 (.A1(n_5_183), .A2(n_5_3895), .ZN(n_5_3897));
   INV_X1 i_5_4747 (.A(n_5_3897), .ZN(n_5_3899));
   NAND3_X1 i_5_4420 (.A1(n_5_4628), .A2(n_5_4625), .A3(n_5_3899), .ZN(n_5_3911));
   NAND2_X1 i_5_4622 (.A1(n_5_132), .A2(n_5_125), .ZN(n_5_3912));
   INV_X1 i_5_4623 (.A(n_5_3912), .ZN(n_5_3913));
   NAND3_X1 i_5_4624 (.A1(n_5_526), .A2(n_5_347), .A3(n_5_3913), .ZN(n_5_3914));
   INV_X1 i_5_4669 (.A(m[14]), .ZN(n_5_3922));
   XNOR2_X1 i_5_4715 (.A(n_5_464), .B(n_5_3922), .ZN(n_5_3923));
   XNOR2_X1 i_5_4745 (.A(n_5_461), .B(n_5_3923), .ZN(n_5_3925));
   XNOR2_X1 i_5_160 (.A(n_5_3947), .B(m[8]), .ZN(n_5_3945));
   NOR2_X1 i_5_4272 (.A1(n_5_3947), .A2(n_60), .ZN(n_5_3956));
   NAND2_X1 i_5_4519 (.A1(n_5_4751), .A2(n_5_218), .ZN(n_5_3960));
   NAND3_X1 i_5_4636 (.A1(n_5_462), .A2(n_5_456), .A3(n_5_460), .ZN(n_5_3983));
   NAND3_X1 i_5_4733 (.A1(n_5_462), .A2(n_5_456), .A3(n_5_460), .ZN(n_5_3984));
   NAND2_X1 i_5_4293 (.A1(n_5_3984), .A2(n_76), .ZN(n_5_3985));
   OAI22_X1 i_5_1093 (.A1(n_5_81), .A2(n_5_28), .B1(n_5_82), .B2(n_5_130), 
      .ZN(n_5_3857));
   NAND2_X1 i_5_4639 (.A1(n_5_3930), .A2(n_69), .ZN(n_5_3997));
   OAI21_X1 i_5_4663 (.A(n_5_310), .B1(n_5_4792), .B2(n_5_4753), .ZN(n_5_4008));
   INV_X1 i_5_4675 (.A(n_5_3911), .ZN(n_5_4009));
   NAND2_X1 i_5_4226 (.A1(n_5_3930), .A2(n_69), .ZN(n_5_4055));
   NAND2_X1 i_5_4294 (.A1(n_5_3911), .A2(n_5_310), .ZN(n_5_4058));
   OAI21_X1 i_5_4453 (.A(n_5_4055), .B1(n_5_4058), .B2(n_5_4795), .ZN(n_5_4231));
   NAND2_X1 i_5_4501 (.A1(n_5_336), .A2(n_5_4231), .ZN(n_5_4247));
   XNOR2_X1 i_5_4505 (.A(n_5_334), .B(n_5_4231), .ZN(n_5_4255));
   OAI21_X1 i_5_4538 (.A(n_5_4247), .B1(n_5_4255), .B2(n_5_336), .ZN(n_5_4258));
   XNOR2_X1 i_5_4692 (.A(n_5_364), .B(n_5_716), .ZN(n_5_4261));
   XNOR2_X1 i_5_4677 (.A(n_5_364), .B(n_5_716), .ZN(n_5_4267));
   NAND2_X1 i_5_4680 (.A1(n_5_4267), .A2(n_5_197), .ZN(n_5_4268));
   NAND2_X1 i_5_4454 (.A1(n_5_702), .A2(m[6]), .ZN(n_5_4291));
   NAND2_X1 i_5_4562 (.A1(n_5_122), .A2(n_5_126), .ZN(n_5_4298));
   INV_X1 i_5_4429 (.A(n_5_711), .ZN(n_5_4301));
   INV_X1 i_5_4732 (.A(m[6]), .ZN(n_5_4354));
   NAND2_X1 i_5_4475 (.A1(n_5_4301), .A2(n_5_4354), .ZN(n_5_4362));
   NAND2_X1 i_5_4573 (.A1(n_5_419), .A2(n_55), .ZN(n_5_4363));
   INV_X1 i_5_4600 (.A(n_5_739), .ZN(n_5_4369));
   OAI21_X1 i_5_4602 (.A(n_5_728), .B1(n_5_419), .B2(n_55), .ZN(n_5_4370));
   OAI21_X1 i_5_4627 (.A(n_5_4363), .B1(n_5_4369), .B2(n_5_4370), .ZN(n_5_4371));
   NAND2_X1 i_5_4681 (.A1(n_5_3891), .A2(n_5_3946), .ZN(n_5_4380));
   INV_X1 i_5_4349 (.A(n_5_4380), .ZN(n_5_4381));
   INV_X1 i_5_4513 (.A(n_5_43), .ZN(n_5_4382));
   NAND2_X1 i_5_4679 (.A1(n_5_4727), .A2(m[0]), .ZN(n_5_4390));
   INV_X1 i_5_218 (.A(n_5_218), .ZN(n_5_4391));
   INV_X1 i_5_230 (.A(n_5_250), .ZN(n_5_4405));
   NAND2_X1 i_5_271 (.A1(n_5_226), .A2(n_5_252), .ZN(n_5_4409));
   AOI21_X1 i_5_4462 (.A(n_5_4391), .B1(n_5_4405), .B2(n_5_4409), .ZN(n_5_4410));
   INV_X1 i_5_3850 (.A(n_5_217), .ZN(n_5_4411));
   NAND2_X1 i_5_4463 (.A1(n_5_4747), .A2(n_5_4411), .ZN(n_5_4418));
   INV_X1 i_5_4762 (.A(n_5_197), .ZN(n_5_4419));
   NAND2_X1 i_5_4464 (.A1(n_5_4411), .A2(n_5_4419), .ZN(n_5_4420));
   AOI22_X1 i_5_34 (.A1(n_5_531), .A2(n_5_4410), .B1(n_5_4418), .B2(n_5_4420), 
      .ZN(n_5_4421));
   NAND3_X1 i_5_4333 (.A1(n_5_363), .A2(n_5_524), .A3(n_5_136), .ZN(n_5_4439));
   XNOR2_X1 i_5_4378 (.A(n_5_4439), .B(m[10]), .ZN(n_5_4485));
   XNOR2_X1 i_5_4382 (.A(n_5_4439), .B(n_73), .ZN(n_5_3931));
   NAND3_X1 i_5_4396 (.A1(n_5_363), .A2(n_5_524), .A3(n_5_136), .ZN(n_5_4509));
   NAND2_X1 i_5_4068 (.A1(n_5_381), .A2(n_5_242), .ZN(n_5_4532));
   NAND2_X1 i_5_4757 (.A1(n_5_243), .A2(m[14]), .ZN(n_5_4535));
   INV_X1 i_5_4587 (.A(n_5_263), .ZN(n_5_4536));
   AOI22_X1 i_5_4640 (.A1(n_5_243), .A2(m[14]), .B1(n_5_381), .B2(n_5_242), 
      .ZN(n_5_4537));
   NAND2_X1 i_5_4758 (.A1(n_5_4536), .A2(n_5_4537), .ZN(n_5_4539));
   NAND3_X1 i_5_4482 (.A1(n_5_4362), .A2(n_5_122), .A3(n_5_126), .ZN(n_5_3932));
   NAND2_X1 i_5_4483 (.A1(n_5_702), .A2(m[6]), .ZN(n_5_3935));
   NAND3_X1 i_5_4492 (.A1(n_5_546), .A2(n_5_4540), .A3(n_5_578), .ZN(n_5_4543));
   XNOR2_X1 i_5_4506 (.A(n_5_4543), .B(m[7]), .ZN(n_5_3936));
   NOR2_X1 i_5_4402 (.A1(n_5_4543), .A2(n_69), .ZN(n_5_4551));
   XNOR2_X1 i_5_4523 (.A(n_5_4543), .B(n_69), .ZN(n_5_4552));
   NOR2_X1 i_5_4339 (.A1(n_5_3961), .A2(m[7]), .ZN(n_5_3858));
   NAND3_X1 i_5_4524 (.A1(n_5_546), .A2(n_5_4540), .A3(n_5_578), .ZN(n_5_3961));
   XNOR2_X1 i_5_4697 (.A(n_5_455), .B(n_5_626), .ZN(n_5_4557));
   NAND2_X1 i_5_4698 (.A1(n_5_4557), .A2(n_5_378), .ZN(n_5_4558));
   NAND2_X1 i_5_4419 (.A1(n_5_4665), .A2(m[10]), .ZN(n_5_4576));
   INV_X1 i_5_4435 (.A(n_5_539), .ZN(n_5_4578));
   NOR2_X1 i_5_4449 (.A1(n_5_175), .A2(n_5_176), .ZN(n_5_4590));
   OAI21_X1 i_5_4759 (.A(n_5_4576), .B1(n_5_4578), .B2(n_5_4590), .ZN(n_5_4597));
   INV_X1 i_5_4511 (.A(n_5_353), .ZN(n_5_4602));
   NAND2_X1 i_5_4049 (.A1(n_5_646), .A2(n_5_188), .ZN(n_5_3859));
   NAND2_X1 i_5_4676 (.A1(n_5_60), .A2(n_5_79), .ZN(n_5_4609));
   NAND3_X1 i_5_4090 (.A1(n_5_4525), .A2(n_5_4800), .A3(n_5_625), .ZN(n_5_4610));
   NAND2_X1 i_5_4695 (.A1(n_5_4382), .A2(n_5_4390), .ZN(n_5_4617));
   NAND2_X1 i_5_4391 (.A1(n_5_4382), .A2(n_5_4390), .ZN(n_5_4618));
   NAND2_X1 i_5_4392 (.A1(n_5_60), .A2(n_5_79), .ZN(n_5_4619));
   NAND3_X1 i_5_4397 (.A1(n_5_4525), .A2(n_5_4800), .A3(n_5_625), .ZN(n_5_4623));
   NAND3_X1 i_5_4425 (.A1(n_5_4618), .A2(n_5_4619), .A3(n_5_4623), .ZN(n_5_3860));
   NAND2_X1 i_5_4543 (.A1(n_5_377), .A2(n_5_197), .ZN(n_5_4625));
   NAND2_X1 i_5_4580 (.A1(n_5_261), .A2(n_5_218), .ZN(n_5_4628));
   NAND2_X1 i_5_4582 (.A1(n_5_377), .A2(n_5_197), .ZN(n_5_4629));
   NAND2_X1 i_5_4583 (.A1(n_5_261), .A2(n_5_218), .ZN(n_5_4630));
   NAND3_X1 i_5_4584 (.A1(n_5_4629), .A2(n_5_4630), .A3(n_5_183), .ZN(n_5_4638));
   NAND3_X1 i_5_4444 (.A1(n_5_701), .A2(n_5_4268), .A3(n_5_184), .ZN(n_5_4643));
   INV_X1 i_5_4473 (.A(n_5_4643), .ZN(n_5_4650));
   NAND2_X1 i_5_4634 (.A1(n_5_4643), .A2(m[8]), .ZN(n_5_4651));
   NAND2_X1 i_5_4688 (.A1(n_5_4643), .A2(n_60), .ZN(n_5_4652));
   NAND3_X1 i_5_4770 (.A1(n_5_701), .A2(n_5_4268), .A3(n_5_184), .ZN(n_5_4660));
   NAND2_X1 i_5_4451 (.A1(n_5_249), .A2(n_5_252), .ZN(n_5_4661));
   NAND2_X1 i_5_4495 (.A1(n_5_4532), .A2(n_5_4535), .ZN(n_5_4662));
   NAND2_X1 i_5_4510 (.A1(n_5_4661), .A2(n_5_4662), .ZN(n_5_4664));
   NAND3_X1 i_5_4386 (.A1(n_5_3960), .A2(n_5_3959), .A3(n_5_196), .ZN(n_5_4665));
   NAND3_X1 i_5_4641 (.A1(n_5_3960), .A2(n_5_3959), .A3(n_5_196), .ZN(n_5_4666));
   INV_X1 i_5_4666 (.A(n_5_4666), .ZN(n_5_4667));
   NAND2_X1 i_5_4385 (.A1(n_5_439), .A2(n_5_440), .ZN(n_5_4668));
   OR2_X1 i_5_4390 (.A1(m[11]), .A2(n_5_293), .ZN(n_5_4691));
   INV_X1 i_5_4428 (.A(m[11]), .ZN(n_5_4692));
   NOR2_X1 i_5_4437 (.A1(n_5_440), .A2(n_5_4692), .ZN(n_5_4693));
   NAND2_X1 i_5_4497 (.A1(n_5_440), .A2(n_5_4692), .ZN(n_5_4708));
   AOI21_X1 i_5_4771 (.A(n_5_4693), .B1(n_5_293), .B2(n_5_4708), .ZN(n_5_4716));
   NOR2_X1 i_5_4772 (.A1(n_5_293), .A2(m[11]), .ZN(n_5_4717));
   OAI21_X1 i_5_4773 (.A(n_5_4716), .B1(n_5_439), .B2(n_5_4717), .ZN(n_5_4719));
   NAND2_X1 i_5_4761 (.A1(n_5_4539), .A2(n_5_4664), .ZN(n_5_4722));
   OAI21_X1 i_5_4704 (.A(n_5_325), .B1(n_5_326), .B2(n_5_525), .ZN(n_5_4723));
   NAND2_X1 i_5_4426 (.A1(n_5_4723), .A2(n_5_95), .ZN(n_5_3861));
   INV_X1 i_5_4642 (.A(n_5_197), .ZN(n_5_4725));
   NOR2_X1 i_5_4737 (.A1(n_5_374), .A2(n_5_4725), .ZN(n_5_4736));
   OAI21_X1 i_5_4763 (.A(n_5_221), .B1(n_5_373), .B2(n_5_4725), .ZN(n_5_4737));
   NOR2_X1 i_5_4768 (.A1(n_5_4736), .A2(n_5_4737), .ZN(n_5_4738));
   INV_X1 i_5_4769 (.A(n_5_218), .ZN(n_5_4739));
   OAI21_X1 i_5_4774 (.A(n_5_4738), .B1(n_5_4722), .B2(n_5_4739), .ZN(n_5_4740));
   NAND2_X1 i_5_4591 (.A1(n_5_4801), .A2(n_5_14), .ZN(n_5_4741));
   NAND2_X1 i_5_4635 (.A1(n_5_27), .A2(n_5_15), .ZN(n_5_4742));
   NAND3_X1 i_5_4652 (.A1(n_5_4741), .A2(n_5_4742), .A3(n_5_22), .ZN(n_90));
   NAND2_X1 i_5_4409 (.A1(n_5_29), .A2(n_5_15), .ZN(n_5_4743));
   INV_X1 i_5_326 (.A(n_5_24), .ZN(n_5_4744));
   AOI21_X1 i_5_4303 (.A(n_5_4744), .B1(n_5_117), .B2(n_5_14), .ZN(n_5_4745));
   NAND2_X1 i_5_4648 (.A1(n_5_4743), .A2(n_5_4745), .ZN(n_91));
   INV_X1 i_5_4504 (.A(n_5_579), .ZN(n_5_4746));
   XNOR2_X1 i_5_4752 (.A(n_5_4746), .B(n_5_581), .ZN(n_5_4747));
   NAND3_X1 i_5_4411 (.A1(n_5_3531), .A2(n_5_185), .A3(n_5_192), .ZN(n_5_4748));
   NAND3_X1 i_5_4601 (.A1(n_5_3531), .A2(n_5_185), .A3(n_5_192), .ZN(n_5_4749));
   INV_X1 i_5_4776 (.A(n_5_4749), .ZN(n_5_4750));
   XNOR2_X1 i_5_601 (.A(n_5_528), .B(n_5_225), .ZN(n_5_4751));
   XNOR2_X1 i_5_4440 (.A(n_5_225), .B(n_5_528), .ZN(n_5_4752));
   NAND2_X1 i_5_4450 (.A1(n_5_4752), .A2(n_5_218), .ZN(n_5_878));
   INV_X1 i_5_4707 (.A(n_5_100), .ZN(n_5_4754));
   XNOR2_X1 i_5_4720 (.A(n_5_4298), .B(n_5_4754), .ZN(n_5_4755));
   NAND2_X1 i_5_4721 (.A1(n_5_4755), .A2(n_5_14), .ZN(n_5_4756));
   NAND3_X1 i_5_4596 (.A1(n_5_418), .A2(n_5_452), .A3(n_5_410), .ZN(n_5_4757));
   XNOR2_X1 i_5_4626 (.A(n_5_4757), .B(m[8]), .ZN(n_5_4758));
   OR2_X1 i_5_4572 (.A1(n_5_4757), .A2(m[8]), .ZN(n_5_4759));
   NAND2_X1 i_5_4646 (.A1(n_5_4757), .A2(m[8]), .ZN(n_5_4760));
   AOI21_X1 i_5_4647 (.A(n_5_376), .B1(n_5_4757), .B2(n_5_375), .ZN(n_5_4761));
   NAND3_X1 i_5_4779 (.A1(n_5_418), .A2(n_5_452), .A3(n_5_410), .ZN(n_5_4762));
   NAND3_X1 i_5_4590 (.A1(n_5_163), .A2(n_5_162), .A3(n_5_181), .ZN(n_5_4763));
   INV_X1 i_5_4594 (.A(n_5_4037), .ZN(n_5_4764));
   INV_X1 i_5_4630 (.A(n_5_182), .ZN(n_5_4765));
   NAND3_X1 i_5_4643 (.A1(n_5_163), .A2(n_5_162), .A3(n_5_181), .ZN(n_5_4766));
   INV_X1 i_5_4780 (.A(n_5_4037), .ZN(n_5_4767));
   INV_X1 i_5_4781 (.A(n_5_182), .ZN(n_5_4768));
   NAND2_X1 i_5_4509 (.A1(n_5_157), .A2(n_5_158), .ZN(n_5_4259));
   INV_X1 i_5_4539 (.A(n_5_4037), .ZN(n_5_4260));
   NAND2_X1 i_5_4588 (.A1(n_5_157), .A2(n_5_158), .ZN(n_5_4279));
   INV_X1 i_5_4777 (.A(n_5_182), .ZN(n_5_4320));
   NAND2_X1 i_5_4581 (.A1(n_5_700), .A2(n_5_420), .ZN(n_5_4774));
   NAND2_X1 i_5_4595 (.A1(n_5_438), .A2(n_5_378), .ZN(n_5_4775));
   NAND2_X1 i_5_4644 (.A1(n_5_700), .A2(n_5_420), .ZN(n_5_4776));
   NAND2_X1 i_5_4645 (.A1(n_5_438), .A2(n_5_378), .ZN(n_5_4777));
   NAND3_X1 i_5_4709 (.A1(n_5_4776), .A2(n_5_4777), .A3(n_5_515), .ZN(n_5_4778));
   INV_X1 i_5_4342 (.A(n_5_684), .ZN(n_5_4779));
   AOI21_X1 i_5_4359 (.A(n_5_4766), .B1(n_5_4767), .B2(n_5_4768), .ZN(n_5_4780));
   INV_X1 i_5_4376 (.A(n_5_692), .ZN(n_5_4781));
   INV_X1 i_5_4417 (.A(n_5_684), .ZN(n_5_4782));
   AOI21_X1 i_5_4786 (.A(n_5_4766), .B1(n_5_4767), .B2(n_5_4768), .ZN(n_5_4783));
   INV_X1 i_5_4787 (.A(n_5_692), .ZN(n_5_4784));
   OAI21_X1 i_5_4788 (.A(n_5_4782), .B1(n_5_4783), .B2(n_5_4784), .ZN(n_5_4785));
   NAND2_X1 i_5_4104 (.A1(n_5_498), .A2(n_5_436), .ZN(n_5_4786));
   INV_X1 i_5_4105 (.A(n_5_4786), .ZN(n_5_4787));
   XNOR2_X1 i_5_4331 (.A(n_5_532), .B(n_5_265), .ZN(n_5_4788));
   NAND2_X1 i_5_4520 (.A1(n_5_4788), .A2(n_5_188), .ZN(n_5_4789));
   NAND2_X1 i_5_4503 (.A1(n_5_294), .A2(n_5_177), .ZN(n_5_619));
   NAND2_X1 i_5_4612 (.A1(n_5_294), .A2(n_5_177), .ZN(n_5_843));
   OAI21_X1 i_5_4678 (.A(n_5_232), .B1(n_5_429), .B2(n_5_270), .ZN(n_5_3937));
   NAND2_X1 i_5_4789 (.A1(n_5_843), .A2(n_5_3937), .ZN(n_5_4037));
   XNOR2_X1 i_5_4518 (.A(n_5_4608), .B(n_5_201), .ZN(n_5_4040));
   NAND2_X1 i_5_4427 (.A1(n_5_4605), .A2(n_5_95), .ZN(n_5_4525));
   OR2_X1 i_5_4742 (.A1(n_5_293), .A2(n_76), .ZN(n_5_4579));
   NAND2_X1 i_5_4748 (.A1(n_5_293), .A2(n_76), .ZN(n_5_4790));
   XNOR2_X1 i_5_4778 (.A(n_5_293), .B(n_76), .ZN(n_5_4791));
   NAND2_X1 i_5_4750 (.A1(n_5_842), .A2(n_5_387), .ZN(n_5_3771));
   NAND2_X1 i_5_4751 (.A1(n_5_421), .A2(n_5_602), .ZN(n_5_3839));
   NAND2_X1 i_5_4753 (.A1(n_5_3771), .A2(n_5_3839), .ZN(n_5_3840));
   NAND2_X1 i_5_4713 (.A1(n_5_367), .A2(n_5_197), .ZN(n_5_3841));
   NAND2_X1 i_5_4724 (.A1(n_5_367), .A2(n_5_197), .ZN(n_5_3959));
   NAND3_X1 i_5_4725 (.A1(n_5_3841), .A2(n_5_878), .A3(n_5_196), .ZN(n_5_3982));
   XNOR2_X1 i_5_4749 (.A(n_5_876), .B(n_5_873), .ZN(n_5_4222));
   XNOR2_X1 i_5_4760 (.A(n_5_873), .B(n_5_876), .ZN(n_5_4447));
   NAND2_X1 i_5_4791 (.A1(n_5_4447), .A2(n_5_378), .ZN(n_5_4600));
   NAND2_X1 i_5_4608 (.A1(n_5_37), .A2(n_5_15), .ZN(n_5_4613));
   NAND2_X1 i_5_4754 (.A1(n_5_38), .A2(n_5_14), .ZN(n_5_4654));
   NAND3_X1 i_5_4755 (.A1(n_5_4613), .A2(n_5_4654), .A3(n_5_25), .ZN(n_92));
   BUF_X1 rt_shieldBuf__2__2__22 (.A(n_56), .Z(n_5_4701));
   NOR2_X1 i_5_4144 (.A1(n_5_323), .A2(n_5_346), .ZN(n_5_4753));
   NAND2_X1 i_5_4158 (.A1(n_5_285), .A2(n_5_365), .ZN(n_5_4792));
   NOR2_X1 i_5_4360 (.A1(n_5_323), .A2(n_5_346), .ZN(n_5_4793));
   NAND2_X1 i_5_4792 (.A1(n_5_285), .A2(n_5_365), .ZN(n_5_4794));
   NOR2_X1 i_5_4793 (.A1(n_5_4793), .A2(n_5_4794), .ZN(n_5_4795));
   INV_X1 i_5_4726 (.A(n_5_496), .ZN(n_5_4326));
   NAND3_X1 i_5_4730 (.A1(n_5_156), .A2(n_5_174), .A3(n_5_239), .ZN(n_5_4327));
   NOR2_X1 i_5_4731 (.A1(n_5_4326), .A2(n_5_4327), .ZN(n_5_4328));
   XNOR2_X1 i_5_4395 (.A(n_5_529), .B(n_5_4603), .ZN(n_5_4494));
   NAND2_X1 i_5_4653 (.A1(n_5_4494), .A2(n_5_188), .ZN(n_5_4540));
   NAND2_X1 i_5_3633 (.A1(n_5_3961), .A2(n_69), .ZN(n_5_4541));
   NAND2_X1 i_5_4683 (.A1(n_5_3961), .A2(n_69), .ZN(n_5_4544));
   INV_X1 i_5_4696 (.A(n_5_4544), .ZN(n_5_4545));
   NOR2_X1 i_5_4783 (.A1(n_5_93), .A2(n_5_4545), .ZN(n_5_4546));
   NAND2_X1 i_5_4358 (.A1(n_5_3930), .A2(m[7]), .ZN(n_5_4547));
   NAND3_X1 i_5_4372 (.A1(n_5_4260), .A2(n_5_4279), .A3(n_5_4320), .ZN(n_5_4550));
   NAND2_X1 i_5_4498 (.A1(n_5_3890), .A2(n_5_4259), .ZN(n_5_4556));
   NAND2_X1 i_5_4507 (.A1(n_5_3930), .A2(m[7]), .ZN(n_5_4599));
   NAND3_X1 i_5_4794 (.A1(n_5_4550), .A2(n_5_4556), .A3(n_5_4599), .ZN(n_5_4603));
   NAND2_X1 i_5_4633 (.A1(n_5_4770), .A2(n_5_188), .ZN(n_5_3891));
   AOI21_X1 i_5_4668 (.A(n_5_576), .B1(n_5_622), .B2(n_5_95), .ZN(n_5_3946));
   AOI21_X1 i_5_4682 (.A(n_5_576), .B1(n_5_622), .B2(n_5_95), .ZN(n_5_4769));
   NAND2_X1 i_5_4714 (.A1(n_5_4802), .A2(n_5_4769), .ZN(n_5_3947));
   XOR2_X1 i_5_4782 (.A(n_5_4726), .B(n_5_3931), .Z(n_5_4772));
   OR2_X1 i_5_4784 (.A1(n_5_4724), .A2(n_5_3706), .ZN(n_5_4773));
   XNOR2_X1 i_5_4565 (.A(n_5_650), .B(n_5_240), .ZN(n_5_4796));
   XNOR2_X1 i_5_4684 (.A(n_5_3873), .B(m[3]), .ZN(n_5_650));
   INV_X1 i_5_4700 (.A(n_5_135), .ZN(n_5_240));
   INV_X1 i_5_4722 (.A(m[3]), .ZN(n_5_4797));
   XNOR2_X1 i_5_4430 (.A(n_5_3873), .B(n_5_4797), .ZN(n_5_4798));
   XNOR2_X1 i_5_4500 (.A(n_5_4798), .B(n_5_135), .ZN(n_5_4799));
   NAND2_X1 i_5_4502 (.A1(n_5_4799), .A2(n_5_188), .ZN(n_5_4800));
   NAND2_X1 i_5_4400 (.A1(n_5_3932), .A2(n_5_3935), .ZN(n_5_4542));
   XNOR2_X1 i_5_4401 (.A(n_5_3936), .B(n_5_4542), .ZN(n_5_4801));
   INV_X1 i_5_4491 (.A(n_5_4803), .ZN(n_5_3955));
   NAND2_X1 i_5_4801 (.A1(n_5_3932), .A2(n_5_3935), .ZN(n_5_4803));
   NAND3_X1 i_5_4521 (.A1(n_5_3859), .A2(n_5_3861), .A3(n_5_180), .ZN(n_5_3966));
   XNOR2_X1 i_5_4522 (.A(n_5_3966), .B(n_58), .ZN(n_5_3974));
   NAND2_X1 i_5_4508 (.A1(n_5_4307), .A2(m[4]), .ZN(n_5_3978));
   XNOR2_X1 i_5_4534 (.A(n_5_3966), .B(m[4]), .ZN(n_5_3995));
   NAND3_X1 i_5_4802 (.A1(n_5_3859), .A2(n_5_3861), .A3(n_5_180), .ZN(n_5_4307));
   XNOR2_X1 i_5_4566 (.A(n_5_87), .B(n_5_3974), .ZN(n_5_4310));
   NAND2_X1 i_5_4571 (.A1(n_5_4310), .A2(n_5_15), .ZN(n_5_4344));
   NAND3_X1 i_5_4603 (.A1(n_5_144), .A2(n_5_210), .A3(n_5_146), .ZN(n_5_4345));
   NAND3_X1 i_5_4656 (.A1(n_5_144), .A2(n_5_210), .A3(n_5_146), .ZN(n_5_4349));
   NAND2_X1 i_5_4699 (.A1(n_5_4349), .A2(m[3]), .ZN(n_5_4372));
   NAND3_X1 i_5_4604 (.A1(n_5_89), .A2(n_5_3860), .A3(n_5_3857), .ZN(n_5_4459));
   INV_X1 i_5_4606 (.A(n_5_4459), .ZN(n_5_4491));
   NAND2_X1 i_5_3657 (.A1(n_5_16), .A2(n_5_15), .ZN(n_5_4502));
   NAND2_X1 i_5_4222 (.A1(n_5_3705), .A2(n_5_14), .ZN(n_5_4521));
   NAND3_X1 i_5_4313 (.A1(n_5_4502), .A2(n_5_4521), .A3(n_5_13), .ZN(n_93));
   NAND2_X1 i_5_4767 (.A1(n_5_3891), .A2(n_5_3946), .ZN(n_5_4523));
   NAND2_X1 i_5_4798 (.A1(n_5_3955), .A2(n_5_96), .ZN(n_5_4555));
   INV_X1 i_5_4799 (.A(n_5_3858), .ZN(n_5_4567));
   INV_X1 i_5_4800 (.A(m[8]), .ZN(n_5_4571));
   NAND3_X1 i_5_4804 (.A1(n_5_3891), .A2(n_5_3946), .A3(n_5_4571), .ZN(n_5_4572));
   NAND3_X1 i_5_4805 (.A1(n_5_4555), .A2(n_5_4567), .A3(n_5_4572), .ZN(n_5_4594));
   OAI22_X1 i_5_4610 (.A1(n_5_316), .A2(n_5_203), .B1(n_5_291), .B2(n_5_209), 
      .ZN(n_5_4604));
   XNOR2_X1 i_5_4613 (.A(n_5_4604), .B(n_5_201), .ZN(n_5_4605));
   OAI22_X1 i_5_4614 (.A1(n_5_316), .A2(n_5_203), .B1(n_5_291), .B2(n_5_209), 
      .ZN(n_5_4608));
   XNOR2_X1 i_5_4654 (.A(n_5_106), .B(n_5_3995), .ZN(n_5_4615));
   NAND2_X1 i_5_4655 (.A1(n_5_4615), .A2(n_5_14), .ZN(n_5_4616));
   NAND2_X1 i_5_4785 (.A1(n_5_3947), .A2(n_60), .ZN(n_5_4624));
   OAI21_X1 i_5_4796 (.A(n_5_26), .B1(n_5_36), .B2(n_5_83), .ZN(n_5_4641));
   OAI21_X1 i_5_4797 (.A(n_5_26), .B1(n_5_36), .B2(n_5_83), .ZN(n_5_4669));
   NAND2_X1 i_5_4807 (.A1(n_5_3947), .A2(n_60), .ZN(n_5_4710));
   NAND2_X1 i_5_4808 (.A1(n_5_4669), .A2(n_5_4710), .ZN(n_5_4720));
   AOI22_X1 i_5_4578 (.A1(n_5_4720), .A2(n_5_88), .B1(n_5_3856), .B2(n_55), 
      .ZN(n_5_4721));
   AOI22_X1 i_5_4703 (.A1(n_5_4720), .A2(n_5_88), .B1(n_5_3856), .B2(n_55), 
      .ZN(n_5_4724));
   OR2_X1 i_5_4766 (.A1(n_5_4721), .A2(n_5_3706), .ZN(n_5_4726));
   NAND3_X1 i_5_4657 (.A1(n_5_127), .A2(n_5_131), .A3(n_5_143), .ZN(n_5_4727));
   NAND3_X1 i_5_4795 (.A1(n_5_131), .A2(n_5_127), .A3(n_5_143), .ZN(n_5_4733));
   NAND2_X1 i_5_4809 (.A1(n_5_4733), .A2(n_5_86), .ZN(n_5_4735));
   XNOR2_X1 i_5_4619 (.A(n_5_465), .B(n_5_189), .ZN(n_5_4770));
   XNOR2_X1 i_5_4625 (.A(n_5_189), .B(n_5_465), .ZN(n_5_4771));
   NAND2_X1 i_5_4810 (.A1(n_5_4771), .A2(n_5_188), .ZN(n_5_4802));
   XNOR2_X1 i_5_4790 (.A(n_5_216), .B(n_5_219), .ZN(n_5_4804));
   XNOR2_X1 i_5_4661 (.A(n_5_216), .B(n_5_219), .ZN(n_5_4805));
   NAND2_X1 i_5_4662 (.A1(n_5_4805), .A2(n_5_197), .ZN(n_5_4806));
   AOI21_X1 i_5_4706 (.A(n_5_123), .B1(n_5_94), .B2(n_5_90), .ZN(n_5_204));
   AOI21_X1 i_5_4685 (.A(n_5_123), .B1(n_5_94), .B2(n_5_90), .ZN(n_5_3862));
   XNOR2_X1 i_5_4756 (.A(n_5_102), .B(n_5_3862), .ZN(n_5_4807));
   OAI21_X1 i_5_4803 (.A(n_5_99), .B1(n_5_211), .B2(n_5_204), .ZN(n_5_4808));
   OAI21_X1 i_5_4811 (.A(n_5_99), .B1(n_5_3862), .B2(n_5_211), .ZN(n_5_4809));
   NAND2_X1 i_5_4764 (.A1(n_5_432), .A2(n_5_443), .ZN(n_5_4810));
   XNOR2_X1 i_5_4765 (.A(n_5_215), .B(n_5_4814), .ZN(n_5_4811));
   NAND3_X1 i_5_4775 (.A1(n_5_4814), .A2(n_5_256), .A3(n_5_199), .ZN(n_5_4812));
   XNOR2_X1 i_5_4806 (.A(n_5_215), .B(n_5_4810), .ZN(n_5_4813));
   NAND2_X1 i_5_4812 (.A1(n_5_432), .A2(n_5_443), .ZN(n_5_4814));
   NAND2_X1 i_7_0 (.A1(n_23), .A2(n_7_20), .ZN(n_7_0));
   NAND2_X1 i_7_1 (.A1(n_7_177), .A2(n_7_23), .ZN(n_7_1));
   NAND2_X1 i_7_2 (.A1(n_7_195), .A2(n_7_27), .ZN(n_7_2));
   NAND3_X1 i_7_3 (.A1(n_7_0), .A2(n_7_1), .A3(n_7_2), .ZN(n_94));
   NAND2_X1 i_7_4 (.A1(n_24), .A2(n_7_20), .ZN(n_7_3));
   NAND2_X1 i_7_5 (.A1(n_7_178), .A2(n_7_23), .ZN(n_7_4));
   NAND2_X1 i_7_6 (.A1(n_15), .A2(n_7_27), .ZN(n_7_5));
   NAND3_X1 i_7_7 (.A1(n_7_3), .A2(n_7_4), .A3(n_7_5), .ZN(n_95));
   NAND2_X1 i_7_8 (.A1(n_25), .A2(n_7_20), .ZN(n_7_6));
   NAND2_X1 i_7_9 (.A1(n_7_179), .A2(n_7_23), .ZN(n_7_7));
   NAND2_X1 i_7_10 (.A1(n_16), .A2(n_7_27), .ZN(n_7_8));
   NAND3_X1 i_7_11 (.A1(n_7_6), .A2(n_7_7), .A3(n_7_8), .ZN(n_96));
   NAND2_X1 i_7_12 (.A1(n_7_180), .A2(n_7_23), .ZN(n_7_9));
   NAND2_X1 i_7_13 (.A1(n_26), .A2(n_7_20), .ZN(n_7_10));
   NAND2_X1 i_7_14 (.A1(n_17), .A2(n_7_27), .ZN(n_7_11));
   NAND3_X1 i_7_15 (.A1(n_7_9), .A2(n_7_10), .A3(n_7_11), .ZN(n_97));
   NAND2_X1 i_7_16 (.A1(n_27), .A2(n_7_20), .ZN(n_7_12));
   NAND2_X1 i_7_17 (.A1(n_7_181), .A2(n_7_23), .ZN(n_7_13));
   NAND2_X1 i_7_18 (.A1(n_18), .A2(n_7_27), .ZN(n_7_14));
   NAND3_X1 i_7_19 (.A1(n_7_12), .A2(n_7_13), .A3(n_7_14), .ZN(n_98));
   NAND2_X1 i_7_20 (.A1(n_28), .A2(n_7_20), .ZN(n_7_15));
   NAND2_X1 i_7_21 (.A1(n_7_185), .A2(n_7_23), .ZN(n_7_16));
   NAND2_X1 i_7_22 (.A1(n_19), .A2(n_7_27), .ZN(n_7_17));
   NAND3_X1 i_7_23 (.A1(n_7_15), .A2(n_7_16), .A3(n_7_17), .ZN(n_99));
   NAND2_X1 i_7_26 (.A1(n_20), .A2(n_7_27), .ZN(n_7_19));
   INV_X1 i_7_28 (.A(r[13]), .ZN(n_7_21));
   NAND2_X1 i_7_29 (.A1(r[14]), .A2(n_7_21), .ZN(n_7_22));
   INV_X1 i_7_30 (.A(n_7_22), .ZN(n_7_20));
   NAND2_X1 i_7_24 (.A1(n_30), .A2(n_7_20), .ZN(n_7_24));
   NOR2_X1 i_7_32 (.A1(r[14]), .A2(n_7_21), .ZN(n_7_23));
   NAND2_X1 i_7_25 (.A1(n_7_182), .A2(n_7_23), .ZN(n_7_26));
   XNOR2_X1 i_7_34 (.A(r[14]), .B(r[13]), .ZN(n_7_27));
   NAND2_X1 i_7_27 (.A1(n_21), .A2(n_7_27), .ZN(n_7_28));
   NAND3_X1 i_7_31 (.A1(n_7_24), .A2(n_7_26), .A3(n_7_28), .ZN(n_100));
   NAND2_X1 i_7_37 (.A1(n_47), .A2(n_89), .ZN(n_7_29));
   INV_X1 i_7_38 (.A(n_7_29), .ZN(result[0]));
   NAND2_X1 i_7_39 (.A1(n_88), .A2(n_47), .ZN(n_7_30));
   INV_X1 i_7_40 (.A(n_7_30), .ZN(result[1]));
   NAND2_X1 i_7_41 (.A1(n_87), .A2(n_47), .ZN(n_7_31));
   INV_X1 i_7_42 (.A(n_7_31), .ZN(result[2]));
   NAND2_X1 i_7_43 (.A1(n_78), .A2(n_47), .ZN(n_7_32));
   INV_X1 i_7_44 (.A(n_7_32), .ZN(result[3]));
   NAND2_X1 i_7_45 (.A1(n_127), .A2(n_47), .ZN(n_7_33));
   INV_X1 i_7_46 (.A(n_7_33), .ZN(result[4]));
   NAND2_X1 i_7_47 (.A1(n_121), .A2(n_47), .ZN(n_7_34));
   INV_X1 i_7_48 (.A(n_7_34), .ZN(result[5]));
   NAND2_X1 i_7_49 (.A1(n_12), .A2(n_47), .ZN(n_7_35));
   INV_X1 i_7_50 (.A(n_7_35), .ZN(result[6]));
   NAND2_X1 i_7_51 (.A1(n_47), .A2(n_7_20), .ZN(n_7_36));
   INV_X1 i_7_52 (.A(n_7_36), .ZN(n_7_37));
   NAND2_X1 i_7_53 (.A1(n_22), .A2(n_7_37), .ZN(n_7_38));
   NAND2_X1 i_7_54 (.A1(n_47), .A2(n_7_23), .ZN(n_7_39));
   INV_X1 i_7_55 (.A(n_7_39), .ZN(n_7_40));
   NAND2_X1 i_7_56 (.A1(n_7_176), .A2(n_7_40), .ZN(n_7_41));
   NAND2_X1 i_7_57 (.A1(n_47), .A2(n_7_27), .ZN(n_7_42));
   INV_X1 i_7_58 (.A(n_7_42), .ZN(n_7_43));
   NAND2_X1 i_7_59 (.A1(n_13), .A2(n_7_43), .ZN(n_7_44));
   NAND3_X1 i_7_60 (.A1(n_7_38), .A2(n_7_41), .A3(n_7_44), .ZN(result[7]));
   NAND2_X1 i_7_61 (.A1(n_23), .A2(n_7_105), .ZN(n_7_45));
   NAND2_X1 i_7_62 (.A1(n_7_177), .A2(n_7_110), .ZN(n_7_46));
   NAND2_X1 i_7_63 (.A1(n_7_195), .A2(n_7_117), .ZN(n_7_47));
   NAND3_X1 i_7_64 (.A1(n_7_45), .A2(n_7_46), .A3(n_7_47), .ZN(n_7_48));
   AOI21_X1 i_7_65 (.A(n_7_48), .B1(n_39), .B2(n_7_95), .ZN(n_7_49));
   INV_X1 i_7_66 (.A(n_31), .ZN(n_7_50));
   OAI21_X1 i_7_67 (.A(n_7_49), .B1(n_7_50), .B2(n_7_99), .ZN(result[8]));
   NAND2_X1 i_7_68 (.A1(n_32), .A2(n_7_100), .ZN(n_7_51));
   NAND2_X1 i_7_69 (.A1(n_40), .A2(n_7_95), .ZN(n_7_52));
   NAND2_X1 i_7_70 (.A1(n_24), .A2(n_7_105), .ZN(n_7_53));
   NAND2_X1 i_7_71 (.A1(n_7_178), .A2(n_7_110), .ZN(n_7_54));
   NAND2_X1 i_7_72 (.A1(n_15), .A2(n_7_117), .ZN(n_7_55));
   NAND3_X1 i_7_73 (.A1(n_7_53), .A2(n_7_54), .A3(n_7_55), .ZN(n_7_56));
   INV_X1 i_7_74 (.A(n_7_56), .ZN(n_7_57));
   NAND3_X1 i_7_75 (.A1(n_7_51), .A2(n_7_52), .A3(n_7_57), .ZN(result[9]));
   NAND2_X1 i_7_76 (.A1(n_33), .A2(n_7_100), .ZN(n_7_58));
   NAND2_X1 i_7_77 (.A1(n_25), .A2(n_7_105), .ZN(n_7_59));
   NAND2_X1 i_7_78 (.A1(n_7_179), .A2(n_7_110), .ZN(n_7_60));
   NAND2_X1 i_7_79 (.A1(n_16), .A2(n_7_117), .ZN(n_7_61));
   NAND3_X1 i_7_80 (.A1(n_7_59), .A2(n_7_60), .A3(n_7_61), .ZN(n_7_62));
   AOI21_X1 i_7_81 (.A(n_7_62), .B1(n_41), .B2(n_7_95), .ZN(n_7_63));
   NAND2_X1 i_7_82 (.A1(n_7_58), .A2(n_7_63), .ZN(result[10]));
   NAND2_X1 i_7_83 (.A1(n_34), .A2(n_7_100), .ZN(n_7_64));
   NAND2_X1 i_7_84 (.A1(n_42), .A2(n_7_95), .ZN(n_7_65));
   NAND2_X1 i_7_85 (.A1(n_26), .A2(n_7_105), .ZN(n_7_66));
   NAND2_X1 i_7_86 (.A1(n_7_180), .A2(n_7_110), .ZN(n_7_67));
   NAND2_X1 i_7_87 (.A1(n_17), .A2(n_7_117), .ZN(n_7_68));
   NAND3_X1 i_7_88 (.A1(n_7_66), .A2(n_7_67), .A3(n_7_68), .ZN(n_7_69));
   INV_X1 i_7_89 (.A(n_7_69), .ZN(n_7_70));
   NAND3_X1 i_7_90 (.A1(n_7_64), .A2(n_7_65), .A3(n_7_70), .ZN(result[11]));
   NAND2_X1 i_7_91 (.A1(n_43), .A2(n_7_95), .ZN(n_7_71));
   NAND2_X1 i_7_92 (.A1(n_35), .A2(n_7_100), .ZN(n_7_72));
   NAND2_X1 i_7_93 (.A1(n_27), .A2(n_7_105), .ZN(n_7_73));
   NAND2_X1 i_7_94 (.A1(n_7_181), .A2(n_7_110), .ZN(n_7_74));
   NAND2_X1 i_7_95 (.A1(n_18), .A2(n_7_117), .ZN(n_7_75));
   NAND3_X1 i_7_96 (.A1(n_7_73), .A2(n_7_74), .A3(n_7_75), .ZN(n_7_76));
   INV_X1 i_7_97 (.A(n_7_76), .ZN(n_7_77));
   NAND3_X1 i_7_98 (.A1(n_7_71), .A2(n_7_72), .A3(n_7_77), .ZN(result[12]));
   NAND2_X1 i_7_99 (.A1(n_44), .A2(n_7_95), .ZN(n_7_78));
   NAND2_X1 i_7_100 (.A1(n_36), .A2(n_7_100), .ZN(n_7_79));
   NAND2_X1 i_7_101 (.A1(n_28), .A2(n_7_105), .ZN(n_7_80));
   NAND2_X1 i_7_102 (.A1(n_7_185), .A2(n_7_110), .ZN(n_7_81));
   NAND2_X1 i_7_103 (.A1(n_19), .A2(n_7_117), .ZN(n_7_82));
   NAND3_X1 i_7_104 (.A1(n_7_80), .A2(n_7_81), .A3(n_7_82), .ZN(n_7_83));
   INV_X1 i_7_105 (.A(n_7_83), .ZN(n_7_84));
   NAND3_X1 i_7_106 (.A1(n_7_78), .A2(n_7_79), .A3(n_7_84), .ZN(result[13]));
   NAND2_X1 i_7_33 (.A1(n_45), .A2(n_7_95), .ZN(n_7_85));
   NAND2_X1 i_7_35 (.A1(n_37), .A2(n_7_100), .ZN(n_7_86));
   NAND2_X1 i_7_36 (.A1(n_7_187), .A2(n_7_110), .ZN(n_7_87));
   NAND2_X1 i_7_110 (.A1(n_29), .A2(n_7_105), .ZN(n_7_88));
   NAND2_X1 i_7_111 (.A1(n_7_194), .A2(n_7_117), .ZN(n_7_89));
   NAND3_X1 i_7_107 (.A1(n_7_87), .A2(n_7_88), .A3(n_7_89), .ZN(n_7_90));
   INV_X1 i_7_108 (.A(n_7_90), .ZN(n_7_91));
   NAND3_X1 i_7_109 (.A1(n_7_85), .A2(n_7_86), .A3(n_7_91), .ZN(result[14]));
   INV_X1 i_7_115 (.A(r[14]), .ZN(n_7_92));
   NOR2_X1 i_7_116 (.A1(r[15]), .A2(n_7_92), .ZN(n_7_93));
   NAND2_X1 i_7_117 (.A1(n_47), .A2(n_7_93), .ZN(n_7_94));
   INV_X1 i_7_118 (.A(n_7_94), .ZN(n_7_95));
   NAND2_X1 i_7_119 (.A1(n_46), .A2(n_7_95), .ZN(n_7_96));
   NAND2_X1 i_7_120 (.A1(r[15]), .A2(n_7_92), .ZN(n_7_97));
   INV_X1 i_7_121 (.A(n_7_97), .ZN(n_7_98));
   NAND2_X1 i_7_122 (.A1(n_47), .A2(n_7_98), .ZN(n_7_99));
   INV_X1 i_7_123 (.A(n_7_99), .ZN(n_7_100));
   NAND2_X1 i_7_124 (.A1(n_38), .A2(n_7_100), .ZN(n_7_101));
   NAND2_X1 i_7_125 (.A1(r[15]), .A2(n_7_20), .ZN(n_7_102));
   INV_X1 i_7_126 (.A(n_7_102), .ZN(n_7_103));
   NAND2_X1 i_7_127 (.A1(n_47), .A2(n_7_103), .ZN(n_7_104));
   INV_X1 i_7_128 (.A(n_7_104), .ZN(n_7_105));
   NAND2_X1 i_7_129 (.A1(n_30), .A2(n_7_105), .ZN(n_7_106));
   NAND2_X1 i_7_130 (.A1(n_7_92), .A2(r[13]), .ZN(n_7_107));
   NOR2_X1 i_7_131 (.A1(r[15]), .A2(n_7_107), .ZN(n_7_108));
   NAND2_X1 i_7_132 (.A1(n_47), .A2(n_7_108), .ZN(n_7_109));
   INV_X1 i_7_133 (.A(n_7_109), .ZN(n_7_110));
   NAND2_X1 i_7_134 (.A1(n_7_182), .A2(n_7_110), .ZN(n_7_111));
   NOR2_X1 i_7_135 (.A1(r[14]), .A2(r[13]), .ZN(n_7_112));
   NAND2_X1 i_7_136 (.A1(r[14]), .A2(r[13]), .ZN(n_7_113));
   INV_X1 i_7_137 (.A(n_7_113), .ZN(n_7_114));
   MUX2_X1 i_7_138 (.A(n_7_112), .B(n_7_114), .S(r[15]), .Z(n_7_115));
   NAND2_X1 i_7_139 (.A1(n_47), .A2(n_7_115), .ZN(n_7_116));
   INV_X1 i_7_140 (.A(n_7_116), .ZN(n_7_117));
   NAND2_X1 i_7_141 (.A1(n_21), .A2(n_7_117), .ZN(n_7_118));
   NAND3_X1 i_7_142 (.A1(n_7_106), .A2(n_7_111), .A3(n_7_118), .ZN(n_7_119));
   INV_X1 i_7_143 (.A(n_7_119), .ZN(n_7_120));
   NAND3_X1 i_7_144 (.A1(n_7_96), .A2(n_7_101), .A3(n_7_120), .ZN(result[15]));
   INV_X1 i_7_145 (.A(n_7_18), .ZN(n_7_176));
   XNOR2_X1 i_7_146 (.A(n_13), .B(m[0]), .ZN(n_7_18));
   XOR2_X1 i_7_147 (.A(n_7_130), .B(n_7_25), .Z(n_7_177));
   NAND2_X1 i_7_148 (.A1(n_7_121), .A2(n_7_131), .ZN(n_7_25));
   INV_X1 i_7_149 (.A(n_7_133), .ZN(n_7_121));
   XNOR2_X1 i_7_150 (.A(n_7_122), .B(n_7_137), .ZN(n_7_178));
   NAND2_X1 i_7_151 (.A1(n_7_156), .A2(n_7_138), .ZN(n_7_122));
   XNOR2_X1 i_7_152 (.A(n_7_123), .B(n_7_129), .ZN(n_7_179));
   NAND2_X1 i_7_153 (.A1(n_7_132), .A2(n_7_148), .ZN(n_7_123));
   XOR2_X1 i_7_154 (.A(n_7_163), .B(n_7_150), .Z(n_7_180));
   XNOR2_X1 i_7_155 (.A(n_7_124), .B(n_7_192), .ZN(n_7_181));
   XNOR2_X1 i_7_156 (.A(n_18), .B(m[5]), .ZN(n_7_124));
   NAND2_X1 i_7_112 (.A1(n_7_169), .A2(n_7_166), .ZN(n_7_182));
   INV_X1 i_7_158 (.A(m[8]), .ZN(n_7_125));
   INV_X1 i_7_113 (.A(n_21), .ZN(n_7_126));
   NAND3_X1 i_7_114 (.A1(n_7_152), .A2(n_7_142), .A3(n_7_128), .ZN(n_7_127));
   OAI21_X1 i_7_157 (.A(n_7_203), .B1(n_19), .B2(m[6]), .ZN(n_7_128));
   AOI21_X1 i_7_164 (.A(n_7_153), .B1(n_7_138), .B2(n_7_143), .ZN(n_7_129));
   NAND2_X1 i_7_168 (.A1(n_13), .A2(m[0]), .ZN(n_7_130));
   NAND2_X1 i_7_169 (.A1(n_14), .A2(m[1]), .ZN(n_7_131));
   NOR2_X1 i_7_170 (.A1(n_14), .A2(m[1]), .ZN(n_7_133));
   NAND2_X1 i_7_171 (.A1(n_15), .A2(m[2]), .ZN(n_7_138));
   OR2_X1 i_7_165 (.A1(n_16), .A2(m[3]), .ZN(n_7_132));
   NAND2_X1 i_7_166 (.A1(n_19), .A2(m[6]), .ZN(n_7_142));
   INV_X1 i_7_167 (.A(n_20), .ZN(n_7_183));
   INV_X1 i_7_177 (.A(m[7]), .ZN(n_7_184));
   INV_X1 i_7_181 (.A(m[6]), .ZN(n_7_144));
   XNOR2_X1 i_7_159 (.A(n_19), .B(n_7_144), .ZN(n_7_145));
   NAND2_X1 i_7_160 (.A1(n_7_145), .A2(n_7_175), .ZN(n_7_146));
   XNOR2_X1 i_7_161 (.A(n_7_162), .B(n_19), .ZN(n_7_147));
   OAI21_X1 i_7_162 (.A(n_7_146), .B1(n_7_147), .B2(n_7_175), .ZN(n_7_185));
   NOR2_X1 i_7_163 (.A1(n_17), .A2(m[4]), .ZN(n_7_135));
   XNOR2_X1 i_7_188 (.A(n_17), .B(m[4]), .ZN(n_7_150));
   NAND2_X1 i_7_173 (.A1(n_7_183), .A2(n_7_184), .ZN(n_7_151));
   NAND2_X1 i_7_190 (.A1(n_20), .A2(m[7]), .ZN(n_7_152));
   NAND2_X1 i_7_180 (.A1(n_7_128), .A2(n_7_142), .ZN(n_7_186));
   NOR2_X1 i_7_196 (.A1(n_15), .A2(m[2]), .ZN(n_7_153));
   INV_X1 i_7_197 (.A(n_15), .ZN(n_7_154));
   INV_X1 i_7_198 (.A(m[2]), .ZN(n_7_155));
   NAND2_X1 i_7_199 (.A1(n_7_154), .A2(n_7_155), .ZN(n_7_156));
   NAND2_X1 i_7_174 (.A1(n_21), .A2(n_7_125), .ZN(n_7_157));
   NAND2_X1 i_7_175 (.A1(n_7_126), .A2(m[8]), .ZN(n_7_158));
   NAND2_X1 i_7_178 (.A1(n_7_126), .A2(m[8]), .ZN(n_7_159));
   NAND2_X1 i_7_179 (.A1(n_21), .A2(n_7_125), .ZN(n_7_160));
   NOR2_X1 i_7_172 (.A1(n_18), .A2(m[5]), .ZN(n_7_161));
   XNOR2_X1 i_7_176 (.A(n_7_161), .B(m[6]), .ZN(n_7_162));
   NAND2_X1 i_7_184 (.A1(n_7_127), .A2(n_7_151), .ZN(n_7_164));
   INV_X1 i_7_185 (.A(n_7_164), .ZN(n_7_165));
   NAND3_X1 i_7_186 (.A1(n_7_158), .A2(n_7_157), .A3(n_7_165), .ZN(n_7_166));
   NAND2_X1 i_7_189 (.A1(n_7_160), .A2(n_7_159), .ZN(n_7_167));
   NAND2_X1 i_7_191 (.A1(n_7_127), .A2(n_7_151), .ZN(n_7_168));
   NAND2_X1 i_7_201 (.A1(n_7_167), .A2(n_7_168), .ZN(n_7_169));
   OAI21_X1 i_7_187 (.A(n_7_170), .B1(n_7_171), .B2(n_7_172), .ZN(n_7_187));
   NAND3_X1 i_7_192 (.A1(n_7_173), .A2(n_7_172), .A3(n_7_174), .ZN(n_7_170));
   AOI22_X1 i_7_193 (.A1(n_7_183), .A2(n_7_184), .B1(n_20), .B2(m[7]), .ZN(
      n_7_171));
   INV_X1 i_7_194 (.A(n_7_186), .ZN(n_7_172));
   NAND2_X1 i_7_195 (.A1(n_7_183), .A2(n_7_184), .ZN(n_7_173));
   NAND2_X1 i_7_204 (.A1(n_7_194), .A2(m[7]), .ZN(n_7_174));
   NAND2_X1 i_7_202 (.A1(n_20), .A2(m[7]), .ZN(n_7_188));
   INV_X1 i_7_203 (.A(n_7_183), .ZN(n_7_189));
   INV_X1 i_7_214 (.A(n_7_184), .ZN(n_7_190));
   OAI21_X1 i_7_207 (.A(n_7_188), .B1(n_7_189), .B2(n_7_190), .ZN(n_7_191));
   XNOR2_X1 i_7_208 (.A(n_7_186), .B(n_7_191), .ZN(n_7_136));
   BUF_X1 rt_shieldBuf__2__2__20 (.A(n_20), .Z(n_7_194));
   BUF_X1 rt_shieldBuf__2__2__21 (.A(n_14), .Z(n_7_195));
   AOI21_X1 i_7_216 (.A(n_7_133), .B1(n_7_131), .B2(n_7_130), .ZN(n_7_137));
   INV_X1 i_7_217 (.A(n_7_133), .ZN(n_7_139));
   NAND2_X1 i_7_218 (.A1(n_7_131), .A2(n_7_130), .ZN(n_7_140));
   NAND2_X1 i_7_219 (.A1(n_7_139), .A2(n_7_140), .ZN(n_7_143));
   NAND2_X1 i_7_213 (.A1(n_16), .A2(m[3]), .ZN(n_7_148));
   NAND2_X1 i_7_209 (.A1(n_16), .A2(m[3]), .ZN(n_7_149));
   INV_X1 i_7_210 (.A(n_7_149), .ZN(n_7_134));
   AOI21_X1 i_7_182 (.A(n_7_192), .B1(n_18), .B2(m[5]), .ZN(n_7_175));
   AOI21_X1 i_7_183 (.A(n_7_135), .B1(n_7_196), .B2(n_7_163), .ZN(n_7_192));
   INV_X1 i_7_200 (.A(n_7_135), .ZN(n_7_193));
   INV_X1 i_7_212 (.A(m[5]), .ZN(n_7_141));
   NOR2_X1 i_7_221 (.A1(n_7_163), .A2(n_7_141), .ZN(n_7_197));
   NOR2_X1 i_7_222 (.A1(n_7_196), .A2(n_7_141), .ZN(n_7_198));
   NAND2_X1 i_7_215 (.A1(n_7_135), .A2(n_7_141), .ZN(n_7_200));
   NAND2_X1 i_7_220 (.A1(n_29), .A2(n_7_20), .ZN(n_7_204));
   NAND2_X1 i_7_223 (.A1(n_7_136), .A2(n_7_23), .ZN(n_7_205));
   NAND3_X1 i_7_224 (.A1(n_7_204), .A2(n_7_205), .A3(n_7_19), .ZN(n_101));
   NAND3_X1 i_7_225 (.A1(n_7_200), .A2(n_7_208), .A3(n_18), .ZN(n_7_201));
   OAI21_X1 i_7_226 (.A(n_7_193), .B1(n_7_197), .B2(n_7_198), .ZN(n_7_202));
   NAND2_X1 i_7_227 (.A1(n_7_201), .A2(n_7_202), .ZN(n_7_203));
   OAI21_X1 i_7_205 (.A(n_7_132), .B1(n_7_134), .B2(n_7_129), .ZN(n_7_163));
   NAND2_X1 i_7_206 (.A1(n_17), .A2(m[4]), .ZN(n_7_196));
   OAI21_X1 i_7_211 (.A(n_7_132), .B1(n_7_134), .B2(n_7_129), .ZN(n_7_199));
   INV_X1 i_7_228 (.A(n_7_141), .ZN(n_7_206));
   AOI21_X1 i_7_229 (.A(n_7_206), .B1(n_17), .B2(m[4]), .ZN(n_7_207));
   NAND2_X1 i_7_230 (.A1(n_7_199), .A2(n_7_207), .ZN(n_7_208));
   INV_X1 i_8_0 (.A(n_8_0), .ZN(n_102));
   XNOR2_X1 i_8_1 (.A(n_125), .B(m[0]), .ZN(n_8_0));
   XNOR2_X1 i_8_2 (.A(n_8_1), .B(n_8_23), .ZN(n_103));
   NAND2_X1 i_8_3 (.A1(n_8_31), .A2(n_8_27), .ZN(n_8_1));
   XNOR2_X1 i_8_4 (.A(n_8_459), .B(n_8_72), .ZN(n_104));
   INV_X1 i_8_5 (.A(m[9]), .ZN(n_8_410));
   NAND2_X1 i_8_6 (.A1(n_8_71), .A2(n_8_36), .ZN(n_8_3));
   NAND2_X1 i_8_7 (.A1(n_8_469), .A2(n_8_20), .ZN(n_8_7));
   NAND2_X1 i_8_8 (.A1(n_8_462), .A2(n_8_21), .ZN(n_8_20));
   AOI21_X1 i_8_9 (.A(n_8_523), .B1(n_8_60), .B2(n_8_86), .ZN(n_8_21));
   INV_X1 i_8_10 (.A(n_8_26), .ZN(n_8_23));
   NAND2_X1 i_8_11 (.A1(n_8_423), .A2(m[0]), .ZN(n_8_26));
   NAND2_X1 i_8_12 (.A1(n_132), .A2(m[8]), .ZN(n_8_36));
   NAND2_X1 i_8_13 (.A1(n_8_82), .A2(n_8_2), .ZN(n_8_8));
   XNOR2_X1 i_8_14 (.A(n_8_39), .B(n_8_8), .ZN(n_105));
   INV_X1 i_8_15 (.A(n_8_514), .ZN(n_8_12));
   NAND2_X1 i_8_17 (.A1(n_8_419), .A2(n_8_88), .ZN(n_8_411));
   INV_X1 i_8_16 (.A(n_8_462), .ZN(n_8_412));
   INV_X1 i_8_21 (.A(n_129), .ZN(n_8_413));
   INV_X1 i_8_22 (.A(m[7]), .ZN(n_8_414));
   NAND2_X1 i_8_24 (.A1(n_8_411), .A2(n_8_415), .ZN(n_8_65));
   NOR2_X1 i_8_26 (.A1(n_8_12), .A2(n_8_538), .ZN(n_8_67));
   OAI21_X1 i_8_27 (.A(n_8_518), .B1(n_8_65), .B2(n_8_67), .ZN(n_106));
   NAND2_X1 i_8_28 (.A1(n_8_480), .A2(m[9]), .ZN(n_8_35));
   INV_X1 i_8_18 (.A(n_123), .ZN(n_8_49));
   INV_X1 i_8_30 (.A(m[1]), .ZN(n_8_54));
   NAND2_X1 i_8_19 (.A1(n_8_49), .A2(n_8_54), .ZN(n_8_31));
   OAI21_X1 i_8_33 (.A(n_8_514), .B1(n_8_53), .B2(n_8_538), .ZN(n_8_70));
   OAI21_X1 i_8_34 (.A(n_8_70), .B1(n_132), .B2(m[8]), .ZN(n_8_71));
   OAI21_X1 i_8_35 (.A(n_8_514), .B1(n_8_53), .B2(n_8_538), .ZN(n_8_72));
   NAND2_X1 i_8_36 (.A1(n_8_35), .A2(n_8_483), .ZN(n_8_76));
   NAND2_X1 i_8_37 (.A1(n_8_76), .A2(n_8_61), .ZN(n_8_77));
   NAND2_X1 i_8_38 (.A1(n_8_480), .A2(m[9]), .ZN(n_8_79));
   NAND3_X1 i_8_39 (.A1(n_8_3), .A2(n_8_79), .A3(n_8_483), .ZN(n_8_80));
   NAND2_X1 i_8_40 (.A1(n_8_77), .A2(n_8_80), .ZN(n_107));
   INV_X1 i_8_41 (.A(n_8_585), .ZN(n_8_415));
   NAND2_X1 i_8_42 (.A1(n_123), .A2(m[1]), .ZN(n_8_27));
   NAND2_X1 i_8_20 (.A1(n_123), .A2(m[1]), .ZN(n_8_28));
   INV_X1 i_8_23 (.A(n_8_28), .ZN(n_8_56));
   OAI21_X1 i_8_45 (.A(n_8_31), .B1(n_8_56), .B2(n_8_23), .ZN(n_8_24));
   XOR2_X1 i_8_46 (.A(n_8_24), .B(n_8_32), .Z(n_108));
   NAND2_X1 i_8_25 (.A1(n_8_25), .A2(n_8_83), .ZN(n_8_82));
   OAI21_X1 i_8_29 (.A(n_8_31), .B1(n_8_56), .B2(n_8_23), .ZN(n_8_83));
   NAND2_X1 i_8_31 (.A1(n_130), .A2(m[4]), .ZN(n_8_416));
   OR2_X1 i_8_32 (.A1(n_122), .A2(m[2]), .ZN(n_8_2));
   NAND2_X1 i_8_43 (.A1(n_122), .A2(m[2]), .ZN(n_8_25));
   XNOR2_X1 i_8_54 (.A(n_122), .B(m[2]), .ZN(n_8_32));
   NOR2_X1 i_8_55 (.A1(n_131), .A2(m[5]), .ZN(n_8_44));
   INV_X1 i_8_56 (.A(n_8_412), .ZN(n_8_46));
   INV_X1 i_8_57 (.A(n_8_44), .ZN(n_8_47));
   NAND2_X1 i_8_58 (.A1(n_8_46), .A2(n_8_47), .ZN(n_8_48));
   NAND2_X1 i_8_59 (.A1(n_8_87), .A2(n_8_48), .ZN(n_8_57));
   NAND2_X1 i_8_60 (.A1(n_8_57), .A2(n_8_75), .ZN(n_109));
   NAND2_X1 i_8_61 (.A1(n_8_469), .A2(n_8_87), .ZN(n_8_417));
   NAND2_X1 i_8_62 (.A1(n_8_469), .A2(n_8_412), .ZN(n_8_418));
   NAND2_X1 i_8_44 (.A1(n_133), .A2(m[6]), .ZN(n_8_419));
   OAI21_X1 i_8_64 (.A(n_8_469), .B1(n_8_412), .B2(n_8_87), .ZN(n_8_88));
   NAND2_X1 i_8_68 (.A1(n_8_585), .A2(n_8_419), .ZN(n_8_43));
   NAND2_X1 i_8_69 (.A1(n_8_7), .A2(n_8_419), .ZN(n_8_45));
   NAND2_X1 i_8_70 (.A1(n_8_43), .A2(n_8_45), .ZN(n_8_53));
   AOI21_X1 i_8_71 (.A(n_8_9), .B1(n_8_8), .B2(n_8_13), .ZN(n_8_58));
   INV_X1 i_8_49 (.A(n_8_60), .ZN(n_8_81));
   XNOR2_X1 i_8_73 (.A(n_8_548), .B(n_8_58), .ZN(n_110));
   AOI21_X1 i_8_52 (.A(n_8_9), .B1(n_8_8), .B2(n_8_13), .ZN(n_8_60));
   INV_X1 i_8_75 (.A(n_8_3), .ZN(n_8_61));
   INV_X1 i_8_76 (.A(m[5]), .ZN(n_8_64));
   XNOR2_X1 i_8_77 (.A(n_131), .B(n_8_64), .ZN(n_8_66));
   OAI21_X1 i_8_78 (.A(n_8_86), .B1(n_8_523), .B2(n_8_60), .ZN(n_8_73));
   NAND2_X1 i_8_79 (.A1(n_8_66), .A2(n_8_73), .ZN(n_8_75));
   INV_X1 i_8_80 (.A(n_8_547), .ZN(n_8_86));
   AOI21_X1 i_8_81 (.A(n_8_547), .B1(n_8_416), .B2(n_8_81), .ZN(n_8_87));
   NAND2_X1 i_8_65 (.A1(n_8_416), .A2(n_8_81), .ZN(n_8_420));
   INV_X1 i_8_66 (.A(n_8_547), .ZN(n_8_421));
   NAND2_X1 i_8_84 (.A1(n_8_577), .A2(n_8_472), .ZN(n_111));
   NOR2_X1 i_8_85 (.A1(n_128), .A2(m[3]), .ZN(n_8_9));
   NAND2_X1 i_8_88 (.A1(n_128), .A2(m[3]), .ZN(n_8_13));
   INV_X1 i_8_93 (.A(m[3]), .ZN(n_8_38));
   XNOR2_X1 i_8_89 (.A(n_128), .B(n_8_38), .ZN(n_8_39));
   INV_X1 i_8_95 (.A(n_8_4), .ZN(n_112));
   OAI21_X1 i_8_96 (.A(n_8_15), .B1(m[0]), .B2(n_125), .ZN(n_8_4));
   XOR2_X1 i_8_97 (.A(n_8_15), .B(n_8_5), .Z(n_113));
   XNOR2_X1 i_8_98 (.A(n_123), .B(n_56), .ZN(n_8_5));
   XOR2_X1 i_8_99 (.A(n_8_11), .B(n_8_580), .Z(n_114));
   NAND2_X1 i_8_100 (.A1(n_8_18), .A2(n_55), .ZN(n_8_17));
   INV_X1 i_8_101 (.A(n_126), .ZN(n_8_18));
   OAI21_X1 i_8_102 (.A(n_8_210), .B1(n_8_40), .B2(n_8_252), .ZN(n_8_11));
   INV_X1 i_8_103 (.A(n_8_457), .ZN(n_8_40));
   NAND2_X1 i_8_104 (.A1(n_8_103), .A2(n_8_98), .ZN(n_115));
   INV_X1 i_8_105 (.A(n_132), .ZN(n_8_19));
   INV_X1 i_8_106 (.A(n_60), .ZN(n_8_6));
   NAND2_X1 i_8_107 (.A1(n_8_41), .A2(n_8_30), .ZN(n_8_10));
   XNOR2_X1 i_8_108 (.A(n_8_10), .B(n_8_34), .ZN(n_116));
   INV_X1 i_8_109 (.A(n_8_545), .ZN(n_8_14));
   BUF_X1 i_8_110 (.A(n_8_16), .Z(n_8_15));
   NAND2_X1 i_8_111 (.A1(n_8_423), .A2(m[0]), .ZN(n_8_16));
   XNOR2_X1 i_8_112 (.A(n_8_105), .B(n_8_22), .ZN(n_117));
   NOR2_X1 i_8_113 (.A1(n_8_37), .A2(n_8_29), .ZN(n_8_22));
   NOR2_X1 i_8_114 (.A1(n_123), .A2(n_56), .ZN(n_8_29));
   OAI21_X1 i_8_115 (.A(n_8_113), .B1(n_8_51), .B2(n_8_109), .ZN(n_118));
   NAND2_X1 i_8_90 (.A1(n_128), .A2(n_65), .ZN(n_8_30));
   NAND2_X1 i_8_117 (.A1(n_8_41), .A2(n_8_34), .ZN(n_8_33));
   OAI21_X1 i_8_118 (.A(n_8_104), .B1(n_8_312), .B2(n_8_37), .ZN(n_8_34));
   AOI22_X1 i_8_119 (.A1(n_123), .A2(n_56), .B1(m[0]), .B2(n_8_423), .ZN(n_8_37));
   OR2_X1 i_8_91 (.A1(n_128), .A2(n_65), .ZN(n_8_41));
   NAND2_X1 i_8_121 (.A1(n_8_91), .A2(n_8_42), .ZN(n_119));
   NAND4_X1 i_8_122 (.A1(n_8_17), .A2(n_8_481), .A3(n_8_92), .A4(n_8_78), 
      .ZN(n_8_42));
   INV_X1 i_8_123 (.A(n_55), .ZN(n_8_422));
   NAND2_X1 i_8_124 (.A1(n_8_33), .A2(n_8_30), .ZN(n_8_63));
   INV_X1 i_8_125 (.A(n_8_63), .ZN(n_8_50));
   AOI21_X1 i_8_126 (.A(n_8_546), .B1(n_8_545), .B2(n_8_50), .ZN(n_8_51));
   OR2_X1 i_8_127 (.A1(n_131), .A2(n_66), .ZN(n_8_52));
   NAND2_X1 i_8_128 (.A1(n_8_50), .A2(n_8_545), .ZN(n_8_182));
   NAND2_X1 i_8_131 (.A1(n_8_33), .A2(n_8_30), .ZN(n_8_55));
   INV_X1 i_8_132 (.A(n_58), .ZN(n_8_59));
   XNOR2_X1 i_8_133 (.A(n_130), .B(n_8_59), .ZN(n_8_62));
   NAND2_X1 i_8_134 (.A1(n_8_33), .A2(n_8_30), .ZN(n_8_68));
   INV_X1 i_8_135 (.A(n_8_68), .ZN(n_8_69));
   NAND2_X1 i_8_137 (.A1(n_129), .A2(n_69), .ZN(n_8_74));
   NAND2_X1 i_8_138 (.A1(n_8_93), .A2(n_8_94), .ZN(n_8_78));
   INV_X1 i_8_139 (.A(n_8_93), .ZN(n_8_84));
   NAND2_X1 i_8_140 (.A1(n_8_19), .A2(n_8_6), .ZN(n_8_85));
   INV_X1 i_8_141 (.A(n_8_94), .ZN(n_8_89));
   AOI22_X1 i_8_142 (.A1(n_8_84), .A2(n_8_85), .B1(n_8_85), .B2(n_8_89), 
      .ZN(n_8_90));
   NAND2_X1 i_8_143 (.A1(n_8_482), .A2(n_8_90), .ZN(n_8_91));
   NAND2_X1 i_8_144 (.A1(n_8_19), .A2(n_8_6), .ZN(n_8_92));
   NAND2_X1 i_8_145 (.A1(n_8_99), .A2(n_8_100), .ZN(n_8_93));
   NAND2_X1 i_8_146 (.A1(n_132), .A2(n_60), .ZN(n_8_94));
   NAND2_X1 i_8_147 (.A1(n_8_19), .A2(n_8_6), .ZN(n_8_95));
   NAND2_X1 i_8_148 (.A1(n_132), .A2(n_60), .ZN(n_8_96));
   NAND2_X1 i_8_149 (.A1(n_8_99), .A2(n_8_100), .ZN(n_8_97));
   NAND3_X1 i_8_150 (.A1(n_8_95), .A2(n_8_96), .A3(n_8_97), .ZN(n_8_98));
   NAND2_X1 i_8_151 (.A1(n_8_11), .A2(n_8_74), .ZN(n_8_99));
   OR2_X1 i_8_152 (.A1(n_129), .A2(n_69), .ZN(n_8_100));
   NOR2_X1 i_8_154 (.A1(n_129), .A2(n_69), .ZN(n_8_101));
   AOI21_X1 i_8_155 (.A(n_8_101), .B1(n_8_11), .B2(n_8_74), .ZN(n_8_102));
   NAND2_X1 i_8_156 (.A1(n_8_571), .A2(n_8_102), .ZN(n_8_103));
   NAND2_X1 i_8_157 (.A1(n_122), .A2(n_59), .ZN(n_8_104));
   XNOR2_X1 i_8_158 (.A(n_122), .B(n_59), .ZN(n_8_105));
   OAI21_X1 i_8_159 (.A(n_8_55), .B1(n_8_14), .B2(n_8_546), .ZN(n_8_106));
   NAND2_X1 i_8_160 (.A1(n_8_69), .A2(n_8_62), .ZN(n_8_107));
   NAND2_X1 i_8_161 (.A1(n_8_106), .A2(n_8_107), .ZN(n_120));
   NOR2_X1 i_8_162 (.A1(n_131), .A2(n_66), .ZN(n_8_108));
   NOR2_X1 i_8_163 (.A1(n_8_108), .A2(n_8_546), .ZN(n_8_183));
   NAND2_X1 i_8_164 (.A1(n_8_52), .A2(n_8_211), .ZN(n_8_109));
   NAND2_X1 i_8_165 (.A1(n_8_50), .A2(n_8_545), .ZN(n_8_110));
   NAND2_X1 i_8_166 (.A1(n_8_211), .A2(n_8_52), .ZN(n_8_111));
   INV_X1 i_8_167 (.A(n_8_546), .ZN(n_8_112));
   NAND3_X1 i_8_168 (.A1(n_8_110), .A2(n_8_111), .A3(n_8_112), .ZN(n_8_113));
   NAND2_X1 i_8_169 (.A1(n_8_128), .A2(n_8_433), .ZN(n_8_114));
   NAND2_X1 i_8_170 (.A1(n_8_484), .A2(n_8_127), .ZN(n_8_115));
   INV_X1 i_8_171 (.A(n_8_115), .ZN(n_8_116));
   AOI21_X1 i_8_172 (.A(n_8_116), .B1(n_8_294), .B2(n_8_434), .ZN(n_8_117));
   NAND2_X1 i_8_173 (.A1(n_8_114), .A2(n_8_117), .ZN(n_121));
   NAND2_X1 i_8_174 (.A1(n_8_134), .A2(n_8_433), .ZN(n_8_118));
   NAND2_X1 i_8_175 (.A1(n_8_295), .A2(n_8_434), .ZN(n_8_119));
   NAND2_X1 i_8_176 (.A1(n_8_485), .A2(n_8_127), .ZN(n_8_120));
   NAND3_X1 i_8_177 (.A1(n_8_118), .A2(n_8_119), .A3(n_8_120), .ZN(n_8_423));
   NAND2_X1 i_8_92 (.A1(n_8_175), .A2(n_8_433), .ZN(n_8_290));
   NAND2_X1 i_8_180 (.A1(n_8_486), .A2(n_8_127), .ZN(n_8_292));
   NAND2_X1 i_8_181 (.A1(n_8_304), .A2(n_8_434), .ZN(n_8_121));
   NAND2_X1 i_8_182 (.A1(n_8_569), .A2(n_8_127), .ZN(n_8_122));
   NAND3_X1 i_8_94 (.A1(n_8_121), .A2(n_8_190), .A3(n_8_122), .ZN(n_122));
   NAND2_X1 i_8_120 (.A1(n_8_513), .A2(n_8_127), .ZN(n_8_424));
   NAND2_X1 i_8_86 (.A1(n_8_302), .A2(n_8_434), .ZN(n_8_425));
   NAND2_X1 i_8_129 (.A1(n_8_493), .A2(n_8_127), .ZN(n_8_123));
   INV_X1 i_8_130 (.A(n_8_123), .ZN(n_8_124));
   AOI21_X1 i_8_188 (.A(n_8_124), .B1(n_8_137), .B2(n_8_433), .ZN(n_8_426));
   NAND2_X1 i_8_194 (.A1(n_8_494), .A2(n_8_127), .ZN(n_8_427));
   NAND2_X1 i_8_196 (.A1(n_8_592), .A2(n_8_127), .ZN(n_8_428));
   NAND2_X1 i_8_47 (.A1(n_8_300), .A2(n_8_434), .ZN(n_8_429));
   NAND2_X1 i_8_48 (.A1(n_8_170), .A2(n_8_433), .ZN(n_8_430));
   NAND2_X1 i_8_199 (.A1(n_8_524), .A2(n_8_127), .ZN(n_8_431));
   NAND2_X1 i_8_116 (.A1(n_8_553), .A2(n_8_127), .ZN(n_8_432));
   INV_X1 i_8_201 (.A(r[11]), .ZN(n_8_125));
   NAND2_X1 i_8_202 (.A1(r[12]), .A2(n_8_125), .ZN(n_8_126));
   INV_X1 i_8_203 (.A(n_8_126), .ZN(n_8_433));
   NOR2_X1 i_8_204 (.A1(r[12]), .A2(n_8_125), .ZN(n_8_434));
   XNOR2_X1 i_8_205 (.A(r[12]), .B(r[11]), .ZN(n_8_127));
   NAND2_X1 i_8_206 (.A1(n_8_504), .A2(n_8_127), .ZN(n_8_435));
   NAND2_X1 i_8_207 (.A1(n_8_298), .A2(n_8_434), .ZN(n_8_436));
   NAND2_X1 i_8_208 (.A1(n_8_145), .A2(n_8_433), .ZN(n_8_437));
   INV_X1 i_8_209 (.A(n_8_129), .ZN(n_8_128));
   XNOR2_X1 i_8_210 (.A(n_8_484), .B(m[0]), .ZN(n_8_129));
   INV_X1 i_8_211 (.A(n_8_196), .ZN(n_8_130));
   NAND2_X1 i_8_153 (.A1(n_8_485), .A2(n_56), .ZN(n_8_131));
   NAND2_X1 i_8_213 (.A1(n_8_130), .A2(n_8_131), .ZN(n_8_132));
   NAND2_X1 i_8_178 (.A1(n_8_484), .A2(m[0]), .ZN(n_8_133));
   XOR2_X1 i_8_215 (.A(n_8_132), .B(n_8_133), .Z(n_8_134));
   AOI21_X1 i_8_179 (.A(n_8_173), .B1(n_8_172), .B2(n_8_176), .ZN(n_8_135));
   XNOR2_X1 i_8_183 (.A(n_8_512), .B(n_8_135), .ZN(n_8_438));
   NAND2_X1 i_8_190 (.A1(n_8_153), .A2(n_8_154), .ZN(n_8_136));
   XNOR2_X1 i_8_191 (.A(n_8_136), .B(n_8_149), .ZN(n_8_137));
   NAND3_X1 i_8_221 (.A1(n_8_165), .A2(n_8_177), .A3(n_8_166), .ZN(n_8_138));
   XNOR2_X1 i_8_195 (.A(n_8_587), .B(n_8_160), .ZN(n_8_439));
   NOR2_X1 i_8_185 (.A1(n_8_553), .A2(n_55), .ZN(n_8_139));
   AOI21_X1 i_8_225 (.A(n_8_139), .B1(n_8_550), .B2(n_8_159), .ZN(n_8_140));
   INV_X1 i_8_226 (.A(n_73), .ZN(n_8_141));
   INV_X1 i_8_227 (.A(n_8_504), .ZN(n_8_142));
   OAI221_X1 i_8_228 (.A(n_8_140), .B1(n_8_504), .B2(n_8_141), .C1(n_73), 
      .C2(n_8_142), .ZN(n_8_143));
   INV_X1 i_8_229 (.A(n_8_140), .ZN(n_8_144));
   NAND2_X1 i_8_230 (.A1(n_8_143), .A2(n_8_186), .ZN(n_8_145));
   NAND2_X1 i_8_184 (.A1(n_8_486), .A2(n_59), .ZN(n_8_192));
   INV_X1 i_8_186 (.A(n_8_192), .ZN(n_8_146));
   NAND2_X1 i_8_50 (.A1(n_8_524), .A2(n_60), .ZN(n_8_147));
   XNOR2_X1 i_8_197 (.A(n_8_524), .B(n_60), .ZN(n_8_148));
   XNOR2_X1 i_8_192 (.A(n_8_493), .B(n_66), .ZN(n_8_149));
   AOI21_X1 i_8_51 (.A(n_8_529), .B1(n_8_147), .B2(n_8_171), .ZN(n_8_150));
   NAND2_X1 i_8_200 (.A1(n_8_139), .A2(n_8_150), .ZN(n_8_151));
   XNOR2_X1 i_8_212 (.A(n_8_550), .B(n_8_150), .ZN(n_8_152));
   NAND2_X1 i_8_242 (.A1(n_8_511), .A2(n_8_135), .ZN(n_8_153));
   NAND2_X1 i_8_243 (.A1(n_8_513), .A2(n_58), .ZN(n_8_154));
   NAND2_X1 i_8_187 (.A1(n_8_135), .A2(n_8_511), .ZN(n_8_155));
   AOI22_X1 i_8_245 (.A1(n_8_493), .A2(n_66), .B1(n_8_513), .B2(n_58), .ZN(
      n_8_156));
   NAND2_X1 i_8_246 (.A1(n_8_171), .A2(n_8_147), .ZN(n_8_157));
   INV_X1 i_8_247 (.A(n_8_529), .ZN(n_8_158));
   NAND2_X1 i_8_248 (.A1(n_8_157), .A2(n_8_158), .ZN(n_8_159));
   NAND2_X1 i_8_222 (.A1(n_8_138), .A2(n_8_188), .ZN(n_8_160));
   NAND2_X1 i_8_87 (.A1(n_8_138), .A2(n_8_188), .ZN(n_8_161));
   INV_X1 i_8_252 (.A(n_8_592), .ZN(n_8_162));
   INV_X1 i_8_253 (.A(n_69), .ZN(n_8_163));
   NAND2_X1 i_8_189 (.A1(n_8_162), .A2(n_8_163), .ZN(n_8_164));
   NAND2_X1 i_8_255 (.A1(n_8_155), .A2(n_8_156), .ZN(n_8_165));
   OR2_X1 i_8_256 (.A1(n_8_493), .A2(n_66), .ZN(n_8_166));
   NOR2_X1 i_8_257 (.A1(n_8_493), .A2(n_66), .ZN(n_8_167));
   INV_X1 i_8_233 (.A(n_8_588), .ZN(n_8_168));
   AOI21_X1 i_8_220 (.A(n_8_168), .B1(n_8_161), .B2(n_8_164), .ZN(n_8_169));
   XOR2_X1 i_8_235 (.A(n_8_148), .B(n_8_169), .Z(n_8_170));
   AOI21_X1 i_8_234 (.A(n_8_168), .B1(n_8_161), .B2(n_8_164), .ZN(n_8_171));
   NAND2_X1 i_8_198 (.A1(n_8_569), .A2(n_65), .ZN(n_8_172));
   NOR2_X1 i_8_214 (.A1(n_8_569), .A2(n_65), .ZN(n_8_173));
   XNOR2_X1 i_8_218 (.A(n_8_569), .B(n_65), .ZN(n_8_174));
   XNOR2_X1 i_8_217 (.A(n_8_198), .B(n_8_194), .ZN(n_8_175));
   INV_X1 i_8_268 (.A(n_8_195), .ZN(n_8_193));
   AOI21_X1 i_8_216 (.A(n_8_146), .B1(n_8_194), .B2(n_8_204), .ZN(n_8_176));
   OR2_X1 i_8_270 (.A1(n_8_494), .A2(n_68), .ZN(n_8_177));
   NOR2_X1 i_8_271 (.A1(n_8_494), .A2(n_68), .ZN(n_8_440));
   NAND2_X1 i_8_272 (.A1(n_8_440), .A2(n_8_199), .ZN(n_8_441));
   INV_X1 i_8_273 (.A(n_8_142), .ZN(n_8_178));
   INV_X1 i_8_274 (.A(n_8_141), .ZN(n_8_179));
   NAND2_X1 i_8_275 (.A1(n_8_178), .A2(n_8_179), .ZN(n_8_180));
   INV_X1 i_8_276 (.A(n_8_504), .ZN(n_8_181));
   INV_X1 i_8_277 (.A(n_73), .ZN(n_8_184));
   NAND2_X1 i_8_278 (.A1(n_8_181), .A2(n_8_184), .ZN(n_8_185));
   NAND3_X1 i_8_279 (.A1(n_8_180), .A2(n_8_144), .A3(n_8_185), .ZN(n_8_186));
   NAND2_X1 i_8_280 (.A1(n_8_494), .A2(n_68), .ZN(n_8_187));
   XNOR2_X1 i_8_281 (.A(n_8_187), .B(n_8_199), .ZN(n_8_442));
   NAND2_X1 i_8_282 (.A1(n_8_494), .A2(n_68), .ZN(n_8_188));
   XNOR2_X1 i_8_219 (.A(n_8_205), .B(n_8_174), .ZN(n_8_189));
   NAND2_X1 i_8_236 (.A1(n_8_189), .A2(n_8_433), .ZN(n_8_190));
   NOR2_X1 i_8_223 (.A1(n_8_485), .A2(n_56), .ZN(n_8_191));
   AOI21_X1 i_8_231 (.A(n_8_191), .B1(n_8_133), .B2(n_8_131), .ZN(n_8_194));
   AOI21_X1 i_8_287 (.A(n_8_191), .B1(n_8_133), .B2(n_8_131), .ZN(n_8_195));
   NOR2_X1 i_8_288 (.A1(n_8_485), .A2(n_56), .ZN(n_8_196));
   NAND2_X1 i_8_238 (.A1(n_8_152), .A2(n_8_151), .ZN(n_8_443));
   INV_X1 i_8_290 (.A(n_8_433), .ZN(n_8_197));
   AOI21_X1 i_8_239 (.A(n_8_197), .B1(n_8_151), .B2(n_8_139), .ZN(n_8_444));
   XNOR2_X1 i_8_232 (.A(n_8_486), .B(n_59), .ZN(n_8_198));
   AOI21_X1 i_8_293 (.A(n_8_167), .B1(n_8_156), .B2(n_8_155), .ZN(n_8_199));
   INV_X1 i_8_294 (.A(n_69), .ZN(n_8_200));
   NAND2_X1 i_8_295 (.A1(n_8_431), .A2(n_8_200), .ZN(n_8_201));
   INV_X1 i_8_296 (.A(n_8_201), .ZN(n_8_445));
   NAND2_X1 i_8_298 (.A1(n_8_182), .A2(n_8_183), .ZN(n_8_202));
   NOR2_X1 i_8_237 (.A1(n_8_486), .A2(n_59), .ZN(n_8_203));
   INV_X1 i_8_240 (.A(n_8_203), .ZN(n_8_204));
   OAI21_X1 i_8_266 (.A(n_8_192), .B1(n_8_193), .B2(n_8_206), .ZN(n_8_205));
   NOR2_X1 i_8_241 (.A1(n_8_486), .A2(n_59), .ZN(n_8_206));
   INV_X1 i_8_305 (.A(n_68), .ZN(n_8_207));
   NAND2_X1 i_8_306 (.A1(n_8_428), .A2(n_8_207), .ZN(n_8_208));
   INV_X1 i_8_307 (.A(n_8_208), .ZN(n_8_209));
   NAND3_X1 i_8_308 (.A1(n_8_539), .A2(n_8_540), .A3(n_8_209), .ZN(n_8_210));
   NAND2_X1 i_8_309 (.A1(n_131), .A2(n_66), .ZN(n_8_211));
   NAND2_X1 i_8_310 (.A1(n_131), .A2(n_66), .ZN(n_8_212));
   INV_X1 i_8_311 (.A(n_8_213), .ZN(n_8_294));
   OAI21_X1 i_8_312 (.A(n_8_222), .B1(m[0]), .B2(n_8_484), .ZN(n_8_213));
   NAND2_X1 i_8_313 (.A1(n_8_493), .A2(m[5]), .ZN(n_8_214));
   NOR2_X1 i_8_314 (.A1(n_8_513), .A2(m[4]), .ZN(n_8_215));
   XOR2_X1 i_8_315 (.A(n_8_222), .B(n_8_216), .Z(n_8_295));
   NAND2_X1 i_8_316 (.A1(n_8_221), .A2(n_8_223), .ZN(n_8_216));
   INV_X1 i_8_317 (.A(n_8_255), .ZN(n_8_217));
   NAND3_X1 i_8_318 (.A1(n_8_267), .A2(n_8_219), .A3(n_8_268), .ZN(n_8_218));
   INV_X1 i_8_319 (.A(n_8_215), .ZN(n_8_219));
   INV_X1 i_8_320 (.A(n_8_241), .ZN(n_8_220));
   INV_X1 i_8_321 (.A(n_8_224), .ZN(n_8_221));
   NAND2_X1 i_8_249 (.A1(n_8_484), .A2(m[0]), .ZN(n_8_222));
   NAND2_X1 i_8_251 (.A1(n_8_485), .A2(m[1]), .ZN(n_8_223));
   NOR2_X1 i_8_267 (.A1(n_8_485), .A2(m[1]), .ZN(n_8_224));
   INV_X1 i_8_289 (.A(n_8_264), .ZN(n_8_225));
   OAI21_X1 i_8_327 (.A(n_8_226), .B1(n_8_237), .B2(n_8_233), .ZN(n_8_298));
   OAI21_X1 i_8_328 (.A(n_8_250), .B1(n_8_260), .B2(n_8_232), .ZN(n_8_226));
   INV_X1 i_8_329 (.A(n_8_241), .ZN(n_8_227));
   OAI21_X1 i_8_254 (.A(n_8_474), .B1(n_8_473), .B2(n_8_229), .ZN(n_8_228));
   NAND2_X1 i_8_260 (.A1(n_8_230), .A2(n_8_246), .ZN(n_8_229));
   NAND3_X1 i_8_261 (.A1(n_8_218), .A2(n_8_214), .A3(n_8_254), .ZN(n_8_230));
   INV_X1 i_8_262 (.A(n_8_591), .ZN(n_8_231));
   NOR2_X1 i_8_335 (.A1(n_8_504), .A2(n_8_234), .ZN(n_8_232));
   NAND2_X1 i_8_336 (.A1(n_8_235), .A2(n_8_258), .ZN(n_8_233));
   INV_X1 i_8_337 (.A(m[10]), .ZN(n_8_234));
   NAND2_X1 i_8_338 (.A1(n_8_236), .A2(m[10]), .ZN(n_8_235));
   INV_X1 i_8_339 (.A(n_8_504), .ZN(n_8_236));
   AOI21_X1 i_8_340 (.A(n_8_238), .B1(n_8_240), .B2(n_8_239), .ZN(n_8_237));
   INV_X1 i_8_341 (.A(n_8_251), .ZN(n_8_238));
   INV_X1 i_8_342 (.A(n_8_220), .ZN(n_8_239));
   INV_X1 i_8_343 (.A(n_8_217), .ZN(n_8_240));
   OAI21_X1 i_8_344 (.A(n_8_242), .B1(n_8_243), .B2(n_8_288), .ZN(n_8_241));
   NAND2_X1 i_8_264 (.A1(n_8_524), .A2(m[8]), .ZN(n_8_242));
   NOR2_X1 i_8_265 (.A1(n_8_524), .A2(m[8]), .ZN(n_8_243));
   XNOR2_X1 i_8_263 (.A(n_8_524), .B(m[8]), .ZN(n_8_244));
   OR2_X1 i_8_193 (.A1(n_8_513), .A2(m[4]), .ZN(n_8_245));
   INV_X1 i_8_330 (.A(n_8_447), .ZN(n_8_246));
   NAND2_X1 i_8_224 (.A1(n_8_493), .A2(m[5]), .ZN(n_8_446));
   NOR2_X1 i_8_323 (.A1(n_8_493), .A2(m[5]), .ZN(n_8_447));
   XNOR2_X1 i_8_324 (.A(n_8_493), .B(m[5]), .ZN(n_8_247));
   NAND2_X1 i_8_356 (.A1(n_8_227), .A2(n_8_251), .ZN(n_8_248));
   NAND2_X1 i_8_357 (.A1(n_8_552), .A2(n_8_251), .ZN(n_8_249));
   NAND2_X1 i_8_358 (.A1(n_8_248), .A2(n_8_249), .ZN(n_8_250));
   NAND2_X1 i_8_334 (.A1(n_8_553), .A2(m[9]), .ZN(n_8_251));
   XNOR2_X1 i_8_353 (.A(n_8_494), .B(m[6]), .ZN(n_8_448));
   XOR2_X1 i_8_331 (.A(n_8_288), .B(n_8_244), .Z(n_8_300));
   NAND2_X1 i_8_363 (.A1(n_8_513), .A2(m[4]), .ZN(n_8_254));
   INV_X1 i_8_364 (.A(n_8_552), .ZN(n_8_255));
   INV_X1 i_8_365 (.A(m[4]), .ZN(n_8_449));
   XNOR2_X1 i_8_244 (.A(n_8_266), .B(n_8_510), .ZN(n_8_450));
   NAND2_X1 i_8_368 (.A1(n_8_504), .A2(n_8_234), .ZN(n_8_258));
   NAND2_X1 i_8_369 (.A1(n_8_504), .A2(n_8_234), .ZN(n_8_259));
   INV_X1 i_8_370 (.A(n_8_259), .ZN(n_8_260));
   NAND2_X1 i_8_325 (.A1(n_8_569), .A2(m[3]), .ZN(n_8_261));
   OR2_X1 i_8_303 (.A1(n_8_486), .A2(m[2]), .ZN(n_8_263));
   NAND2_X1 i_8_269 (.A1(n_8_486), .A2(m[2]), .ZN(n_8_264));
   XNOR2_X1 i_8_283 (.A(n_8_486), .B(m[2]), .ZN(n_8_451));
   NAND2_X1 i_8_284 (.A1(n_8_267), .A2(n_8_268), .ZN(n_8_266));
   NAND2_X1 i_8_377 (.A1(n_8_277), .A2(n_8_261), .ZN(n_8_267));
   OR2_X1 i_8_378 (.A1(n_8_569), .A2(m[3]), .ZN(n_8_268));
   INV_X1 i_8_355 (.A(n_8_261), .ZN(n_8_269));
   INV_X1 i_8_373 (.A(n_8_568), .ZN(n_8_271));
   NAND2_X1 i_8_361 (.A1(n_8_269), .A2(n_8_271), .ZN(n_8_272));
   OAI21_X1 i_8_371 (.A(n_8_272), .B1(n_8_277), .B2(n_8_568), .ZN(n_8_273));
   XOR2_X1 i_8_380 (.A(n_8_247), .B(n_8_274), .Z(n_8_302));
   OAI21_X1 i_8_381 (.A(n_8_245), .B1(n_8_286), .B2(n_8_273), .ZN(n_8_274));
   NAND2_X1 i_8_301 (.A1(n_8_552), .A2(n_8_289), .ZN(n_8_275));
   XNOR2_X1 i_8_302 (.A(n_8_289), .B(n_8_551), .ZN(n_8_276));
   OAI21_X1 i_8_304 (.A(n_8_275), .B1(n_8_276), .B2(n_8_552), .ZN(n_8_452));
   XOR2_X1 i_8_372 (.A(n_8_567), .B(n_8_283), .Z(n_8_304));
   OAI21_X1 i_8_374 (.A(n_8_263), .B1(n_8_225), .B2(n_8_454), .ZN(n_8_277));
   AOI21_X1 i_8_379 (.A(n_8_447), .B1(n_8_455), .B2(n_8_446), .ZN(n_8_453));
   AOI21_X1 i_8_376 (.A(n_8_224), .B1(n_8_223), .B2(n_8_222), .ZN(n_8_281));
   AOI21_X1 i_8_292 (.A(n_8_224), .B1(n_8_223), .B2(n_8_222), .ZN(n_8_454));
   OAI21_X1 i_8_382 (.A(n_8_263), .B1(n_8_225), .B2(n_8_281), .ZN(n_8_283));
   XNOR2_X1 i_8_384 (.A(n_8_513), .B(m[4]), .ZN(n_8_284));
   OAI21_X1 i_8_391 (.A(n_8_245), .B1(n_8_284), .B2(n_8_273), .ZN(n_8_455));
   XNOR2_X1 i_8_385 (.A(n_8_513), .B(m[4]), .ZN(n_8_286));
   AOI21_X1 i_8_332 (.A(n_8_231), .B1(n_8_590), .B2(n_8_228), .ZN(n_8_287));
   AOI21_X1 i_8_333 (.A(n_8_231), .B1(n_8_590), .B2(n_8_228), .ZN(n_8_288));
   OAI21_X1 i_8_346 (.A(n_8_242), .B1(n_8_243), .B2(n_8_287), .ZN(n_8_289));
   XNOR2_X1 i_8_402 (.A(n_8_520), .B(n_8_589), .ZN(n_8_456));
   NAND3_X1 i_8_299 (.A1(n_8_290), .A2(n_8_559), .A3(n_8_292), .ZN(n_123));
   INV_X1 i_8_405 (.A(n_56), .ZN(n_8_308));
   NAND2_X1 i_8_406 (.A1(n_8_292), .A2(n_8_308), .ZN(n_8_309));
   INV_X1 i_8_407 (.A(n_8_309), .ZN(n_8_310));
   NAND3_X1 i_8_408 (.A1(n_8_559), .A2(n_8_290), .A3(n_8_310), .ZN(n_8_311));
   OAI21_X1 i_8_409 (.A(n_8_311), .B1(n_122), .B2(n_59), .ZN(n_8_312));
   NAND2_X1 i_8_410 (.A1(n_8_212), .A2(n_8_202), .ZN(n_8_252));
   NAND2_X1 i_8_411 (.A1(n_8_457), .A2(n_8_210), .ZN(n_8_253));
   NAND2_X1 i_8_412 (.A1(n_8_202), .A2(n_8_212), .ZN(n_8_313));
   XNOR2_X1 i_8_413 (.A(n_8_253), .B(n_8_313), .ZN(n_124));
   NAND2_X1 i_8_418 (.A1(n_8_543), .A2(n_68), .ZN(n_8_457));
   NAND3_X1 i_8_420 (.A1(n_8_554), .A2(n_8_555), .A3(n_8_432), .ZN(n_8_458));
   XNOR2_X1 i_8_421 (.A(n_8_458), .B(m[8]), .ZN(n_8_459));
   NAND3_X1 i_8_347 (.A1(n_8_429), .A2(n_8_430), .A3(n_8_431), .ZN(n_8_460));
   BUF_X1 rt_shieldBuf__2 (.A(n_8_423), .Z(n_125));
   NAND3_X1 i_8_427 (.A1(n_8_561), .A2(n_8_560), .A3(n_8_427), .ZN(n_8_461));
   NAND2_X1 i_8_428 (.A1(n_8_461), .A2(m[5]), .ZN(n_8_462));
   NAND2_X1 i_8_429 (.A1(n_8_442), .A2(n_8_441), .ZN(n_8_463));
   INV_X1 i_8_430 (.A(n_8_433), .ZN(n_8_464));
   AOI21_X1 i_8_431 (.A(n_8_464), .B1(n_8_441), .B2(n_8_440), .ZN(n_8_465));
   INV_X1 i_8_434 (.A(m[5]), .ZN(n_8_466));
   NAND2_X1 i_8_435 (.A1(n_8_427), .A2(n_8_466), .ZN(n_8_467));
   INV_X1 i_8_436 (.A(n_8_467), .ZN(n_8_468));
   NAND3_X1 i_8_437 (.A1(n_8_560), .A2(n_8_561), .A3(n_8_468), .ZN(n_8_469));
   NAND2_X1 i_8_63 (.A1(n_8_415), .A2(n_8_419), .ZN(n_8_470));
   NAND2_X1 i_8_136 (.A1(n_8_417), .A2(n_8_418), .ZN(n_8_471));
   NAND2_X1 i_8_297 (.A1(n_8_470), .A2(n_8_471), .ZN(n_8_472));
   NOR2_X1 i_8_348 (.A1(n_8_494), .A2(m[6]), .ZN(n_8_473));
   NAND2_X1 i_8_349 (.A1(n_8_494), .A2(m[6]), .ZN(n_8_474));
   NAND2_X1 i_8_443 (.A1(n_8_494), .A2(m[6]), .ZN(n_8_475));
   NOR2_X1 i_8_444 (.A1(n_8_494), .A2(m[6]), .ZN(n_8_476));
   OAI21_X1 i_8_445 (.A(n_8_475), .B1(n_8_447), .B2(n_8_476), .ZN(n_8_477));
   NAND3_X1 i_8_446 (.A1(n_8_455), .A2(n_8_475), .A3(n_8_446), .ZN(n_8_478));
   NAND3_X1 i_8_449 (.A1(n_8_436), .A2(n_8_437), .A3(n_8_435), .ZN(n_8_479));
   INV_X1 i_8_450 (.A(n_8_479), .ZN(n_8_480));
   NAND2_X1 i_8_451 (.A1(n_126), .A2(n_8_422), .ZN(n_8_481));
   XNOR2_X1 i_8_452 (.A(n_8_479), .B(n_8_422), .ZN(n_8_482));
   NAND2_X1 i_8_453 (.A1(n_126), .A2(n_8_410), .ZN(n_8_483));
   NAND3_X1 i_8_454 (.A1(n_8_436), .A2(n_8_437), .A3(n_8_435), .ZN(n_126));
   NAND2_X1 i_8_455 (.A1(n_8_405), .A2(n_8_320), .ZN(n_8_256));
   INV_X1 i_8_456 (.A(n_8_256), .ZN(n_8_257));
   AOI21_X1 i_8_457 (.A(n_8_257), .B1(n_0), .B2(n_8_318), .ZN(n_8_262));
   INV_X1 i_8_458 (.A(n_8_262), .ZN(n_8_265));
   AOI21_X1 i_8_459 (.A(n_8_265), .B1(n_8_323), .B2(n_8_315), .ZN(n_8_270));
   INV_X1 i_8_460 (.A(n_8_270), .ZN(n_127));
   NAND2_X1 i_8_461 (.A1(n_1), .A2(n_8_318), .ZN(n_8_278));
   NAND2_X1 i_8_462 (.A1(n_8_325), .A2(n_8_315), .ZN(n_8_279));
   NAND2_X1 i_8_463 (.A1(n_80), .A2(n_8_320), .ZN(n_8_280));
   NAND3_X1 i_8_285 (.A1(n_8_278), .A2(n_8_279), .A3(n_8_280), .ZN(n_8_484));
   NAND2_X1 i_8_465 (.A1(n_8_333), .A2(n_8_315), .ZN(n_8_282));
   NAND2_X1 i_8_466 (.A1(n_2), .A2(n_8_318), .ZN(n_8_285));
   NAND2_X1 i_8_467 (.A1(n_93), .A2(n_8_320), .ZN(n_8_291));
   NAND3_X1 i_8_286 (.A1(n_8_282), .A2(n_8_285), .A3(n_8_291), .ZN(n_8_485));
   NAND2_X1 i_8_291 (.A1(n_3), .A2(n_8_318), .ZN(n_8_293));
   NAND2_X1 i_8_470 (.A1(n_81), .A2(n_8_320), .ZN(n_8_296));
   NAND3_X1 i_8_326 (.A1(n_8_404), .A2(n_8_293), .A3(n_8_296), .ZN(n_8_486));
   NAND2_X1 i_8_351 (.A1(n_4), .A2(n_8_318), .ZN(n_8_487));
   NAND2_X1 i_8_354 (.A1(n_8_334), .A2(n_8_315), .ZN(n_8_488));
   NAND2_X1 i_8_474 (.A1(n_82), .A2(n_8_320), .ZN(n_8_489));
   NAND2_X1 i_8_359 (.A1(n_5), .A2(n_8_318), .ZN(n_8_490));
   NAND2_X1 i_8_360 (.A1(n_8_335), .A2(n_8_315), .ZN(n_8_491));
   NAND2_X1 i_8_478 (.A1(n_83), .A2(n_8_320), .ZN(n_8_492));
   NAND2_X1 i_8_398 (.A1(n_6), .A2(n_8_318), .ZN(n_8_297));
   NAND2_X1 i_8_476 (.A1(n_8_336), .A2(n_8_315), .ZN(n_8_299));
   NAND2_X1 i_8_482 (.A1(n_90), .A2(n_8_320), .ZN(n_8_301));
   NAND3_X1 i_8_477 (.A1(n_8_297), .A2(n_8_299), .A3(n_8_301), .ZN(n_8_493));
   NAND2_X1 i_8_484 (.A1(n_8_337), .A2(n_8_315), .ZN(n_8_303));
   NAND2_X1 i_8_485 (.A1(n_91), .A2(n_8_320), .ZN(n_8_305));
   INV_X1 i_8_486 (.A(n_8_305), .ZN(n_8_306));
   AOI21_X1 i_8_487 (.A(n_8_306), .B1(n_7), .B2(n_8_318), .ZN(n_8_307));
   NAND2_X1 i_8_350 (.A1(n_8_303), .A2(n_8_307), .ZN(n_8_494));
   NAND2_X1 i_8_352 (.A1(n_8), .A2(n_8_318), .ZN(n_8_495));
   NAND2_X1 i_8_362 (.A1(n_8_397), .A2(n_8_315), .ZN(n_8_496));
   NAND2_X1 i_8_491 (.A1(n_84), .A2(n_8_320), .ZN(n_8_497));
   NAND2_X1 i_8_400 (.A1(n_9), .A2(n_8_318), .ZN(n_8_498));
   NAND2_X1 i_8_415 (.A1(n_8_401), .A2(n_8_315), .ZN(n_8_499));
   NAND2_X1 i_8_495 (.A1(n_85), .A2(n_8_320), .ZN(n_8_500));
   NAND2_X1 i_8_387 (.A1(n_8_338), .A2(n_8_315), .ZN(n_8_501));
   NAND2_X1 i_8_388 (.A1(n_10), .A2(n_8_318), .ZN(n_8_502));
   NAND2_X1 i_8_389 (.A1(n_92), .A2(n_8_320), .ZN(n_8_503));
   INV_X1 i_8_501 (.A(r[10]), .ZN(n_8_314));
   NOR2_X1 i_8_502 (.A1(r[11]), .A2(n_8_314), .ZN(n_8_315));
   NAND2_X1 i_8_503 (.A1(n_8_340), .A2(n_8_315), .ZN(n_8_316));
   NAND2_X1 i_8_504 (.A1(r[11]), .A2(n_8_314), .ZN(n_8_317));
   INV_X1 i_8_505 (.A(n_8_317), .ZN(n_8_318));
   NAND2_X1 i_8_506 (.A1(n_11), .A2(n_8_318), .ZN(n_8_319));
   XNOR2_X1 i_8_507 (.A(r[11]), .B(r[10]), .ZN(n_8_320));
   NAND2_X1 i_8_508 (.A1(n_86), .A2(n_8_320), .ZN(n_8_321));
   NAND3_X1 i_8_509 (.A1(n_8_316), .A2(n_8_319), .A3(n_8_321), .ZN(n_8_504));
   BUF_X1 rt_shieldBuf__2__2__23 (.A(n_8_372), .Z(n_8_322));
   INV_X1 i_8_510 (.A(n_8_324), .ZN(n_8_323));
   XNOR2_X1 i_8_511 (.A(n_8_405), .B(m[0]), .ZN(n_8_324));
   XOR2_X1 i_8_512 (.A(n_8_354), .B(n_8_326), .Z(n_8_325));
   NAND2_X1 i_8_513 (.A1(n_8_327), .A2(n_8_355), .ZN(n_8_326));
   INV_X1 i_8_514 (.A(n_8_328), .ZN(n_8_327));
   NOR2_X1 i_8_515 (.A1(n_80), .A2(m[1]), .ZN(n_8_328));
   INV_X1 i_8_516 (.A(m[11]), .ZN(n_8_329));
   INV_X1 i_8_517 (.A(n_86), .ZN(n_8_330));
   NAND2_X1 i_8_518 (.A1(n_86), .A2(n_8_329), .ZN(n_8_331));
   NAND2_X1 i_8_519 (.A1(n_8_330), .A2(m[11]), .ZN(n_8_332));
   XOR2_X1 i_8_520 (.A(n_8_352), .B(n_8_369), .Z(n_8_333));
   INV_X1 i_8_403 (.A(n_8_357), .ZN(n_8_505));
   XNOR2_X1 i_8_395 (.A(n_8_367), .B(n_8_350), .ZN(n_8_334));
   XOR2_X1 i_8_523 (.A(n_8_348), .B(n_8_376), .Z(n_8_335));
   XNOR2_X1 i_8_524 (.A(n_8_395), .B(n_8_347), .ZN(n_8_336));
   XOR2_X1 i_8_525 (.A(n_8_346), .B(n_8_378), .Z(n_8_337));
   XNOR2_X1 i_8_390 (.A(n_8_385), .B(n_8_387), .ZN(n_8_338));
   NAND2_X1 i_8_392 (.A1(n_8_398), .A2(n_8_373), .ZN(n_8_339));
   NAND2_X1 i_8_528 (.A1(n_8_390), .A2(n_8_341), .ZN(n_8_340));
   NAND3_X1 i_8_529 (.A1(n_8_332), .A2(n_8_331), .A3(n_8_407), .ZN(n_8_341));
   NAND2_X1 i_8_530 (.A1(n_8_322), .A2(n_8_343), .ZN(n_8_342));
   NAND2_X1 i_8_531 (.A1(n_8_402), .A2(n_8_398), .ZN(n_8_343));
   INV_X1 i_8_419 (.A(n_8_379), .ZN(n_8_344));
   NAND2_X1 i_8_533 (.A1(n_8_346), .A2(n_8_359), .ZN(n_8_345));
   OAI21_X1 i_8_534 (.A(n_8_393), .B1(n_8_358), .B2(n_8_347), .ZN(n_8_346));
   AOI21_X1 i_8_535 (.A(n_8_364), .B1(n_8_348), .B2(n_8_375), .ZN(n_8_347));
   OAI21_X1 i_8_536 (.A(n_8_365), .B1(n_8_349), .B2(n_8_350), .ZN(n_8_348));
   INV_X1 i_8_537 (.A(n_8_366), .ZN(n_8_349));
   AOI21_X1 i_8_522 (.A(n_8_357), .B1(n_8_371), .B2(n_8_391), .ZN(n_8_350));
   NAND2_X1 i_8_417 (.A1(n_8_352), .A2(n_8_356), .ZN(n_8_351));
   OAI21_X1 i_8_422 (.A(n_8_353), .B1(m[1]), .B2(n_80), .ZN(n_8_352));
   NAND2_X1 i_8_424 (.A1(n_8_355), .A2(n_8_354), .ZN(n_8_353));
   NAND2_X1 i_8_426 (.A1(n_79), .A2(m[0]), .ZN(n_8_354));
   NAND2_X1 i_8_432 (.A1(n_80), .A2(m[1]), .ZN(n_8_355));
   NAND2_X1 i_8_433 (.A1(n_93), .A2(m[2]), .ZN(n_8_356));
   NOR2_X1 i_8_539 (.A1(n_81), .A2(m[3]), .ZN(n_8_357));
   INV_X1 i_8_546 (.A(n_8_394), .ZN(n_8_358));
   NAND2_X1 i_8_547 (.A1(n_91), .A2(m[7]), .ZN(n_8_359));
   OR2_X1 i_8_548 (.A1(n_84), .A2(m[8]), .ZN(n_8_360));
   INV_X1 i_8_549 (.A(m[10]), .ZN(n_8_361));
   INV_X1 i_8_550 (.A(n_8_381), .ZN(n_8_362));
   INV_X1 i_8_551 (.A(n_8_342), .ZN(n_8_363));
   NOR2_X1 i_8_552 (.A1(n_83), .A2(m[5]), .ZN(n_8_364));
   OR2_X1 i_8_553 (.A1(n_82), .A2(m[4]), .ZN(n_8_365));
   NAND2_X1 i_8_554 (.A1(n_82), .A2(m[4]), .ZN(n_8_366));
   XNOR2_X1 i_8_545 (.A(n_82), .B(m[4]), .ZN(n_8_367));
   OR2_X1 i_8_556 (.A1(n_93), .A2(m[2]), .ZN(n_8_368));
   NAND2_X1 i_8_557 (.A1(n_8_368), .A2(n_8_356), .ZN(n_8_369));
   OR2_X1 i_8_438 (.A1(n_93), .A2(m[2]), .ZN(n_8_370));
   NAND2_X1 i_8_558 (.A1(n_8_370), .A2(n_8_351), .ZN(n_8_371));
   OR2_X1 i_8_393 (.A1(n_85), .A2(m[9]), .ZN(n_8_372));
   NAND2_X1 i_8_561 (.A1(n_85), .A2(m[9]), .ZN(n_8_373));
   INV_X1 i_8_562 (.A(m[9]), .ZN(n_8_374));
   NAND2_X1 i_8_563 (.A1(n_83), .A2(m[5]), .ZN(n_8_375));
   XNOR2_X1 i_8_564 (.A(n_83), .B(m[5]), .ZN(n_8_376));
   OR2_X1 i_8_565 (.A1(n_91), .A2(m[7]), .ZN(n_8_377));
   NAND2_X1 i_8_566 (.A1(n_8_380), .A2(n_8_359), .ZN(n_8_378));
   NAND2_X1 i_8_567 (.A1(n_8_377), .A2(n_8_345), .ZN(n_8_379));
   OR2_X1 i_8_568 (.A1(n_91), .A2(m[7]), .ZN(n_8_380));
   NAND2_X1 i_8_569 (.A1(n_92), .A2(m[10]), .ZN(n_8_381));
   INV_X1 i_8_396 (.A(n_92), .ZN(n_8_382));
   INV_X1 i_8_571 (.A(m[10]), .ZN(n_8_383));
   INV_X1 i_8_572 (.A(n_8_361), .ZN(n_8_384));
   OAI22_X1 i_8_397 (.A1(n_8_382), .A2(n_8_383), .B1(n_92), .B2(n_8_384), 
      .ZN(n_8_385));
   NAND2_X1 i_8_439 (.A1(n_8_370), .A2(n_8_351), .ZN(n_8_506));
   NAND2_X1 i_8_399 (.A1(n_8_339), .A2(n_8_372), .ZN(n_8_386));
   INV_X1 i_8_404 (.A(n_8_386), .ZN(n_8_387));
   NAND2_X1 i_8_577 (.A1(n_8_331), .A2(n_8_332), .ZN(n_8_388));
   AOI21_X1 i_8_578 (.A(n_8_362), .B1(n_8_363), .B2(n_8_408), .ZN(n_8_389));
   NAND2_X1 i_8_579 (.A1(n_8_388), .A2(n_8_389), .ZN(n_8_390));
   NAND2_X1 i_8_440 (.A1(n_81), .A2(m[3]), .ZN(n_8_391));
   NAND2_X1 i_8_464 (.A1(n_81), .A2(m[3]), .ZN(n_8_392));
   INV_X1 i_8_468 (.A(n_8_392), .ZN(n_8_507));
   OR2_X1 i_8_583 (.A1(n_90), .A2(m[6]), .ZN(n_8_393));
   NAND2_X1 i_8_584 (.A1(n_90), .A2(m[6]), .ZN(n_8_394));
   XNOR2_X1 i_8_585 (.A(n_90), .B(m[6]), .ZN(n_8_395));
   XNOR2_X1 i_8_586 (.A(n_84), .B(m[8]), .ZN(n_8_396));
   XNOR2_X1 i_8_423 (.A(n_8_399), .B(n_8_344), .ZN(n_8_397));
   OAI21_X1 i_8_588 (.A(n_8_360), .B1(n_8_396), .B2(n_8_344), .ZN(n_8_398));
   XNOR2_X1 i_8_425 (.A(n_84), .B(m[8]), .ZN(n_8_399));
   XNOR2_X1 i_8_590 (.A(n_85), .B(n_8_374), .ZN(n_8_400));
   XNOR2_X1 i_8_591 (.A(n_8_400), .B(n_8_398), .ZN(n_8_401));
   XNOR2_X1 i_8_592 (.A(n_85), .B(n_8_374), .ZN(n_8_402));
   NAND2_X1 i_8_469 (.A1(n_8_351), .A2(n_8_370), .ZN(n_8_403));
   INV_X1 i_8_471 (.A(n_8_403), .ZN(n_8_508));
   NAND2_X1 i_8_366 (.A1(n_8_533), .A2(n_8_315), .ZN(n_8_404));
   BUF_X1 rt_shieldBuf__2__2__18 (.A(n_79), .Z(n_8_405));
   NOR2_X1 i_8_599 (.A1(n_92), .A2(m[10]), .ZN(n_8_406));
   OAI21_X1 i_8_600 (.A(n_8_381), .B1(n_8_342), .B2(n_8_406), .ZN(n_8_407));
   INV_X1 i_8_601 (.A(n_8_409), .ZN(n_8_408));
   NOR2_X1 i_8_602 (.A1(n_92), .A2(m[10]), .ZN(n_8_409));
   NAND3_X1 i_8_367 (.A1(n_8_490), .A2(n_8_491), .A3(n_8_492), .ZN(n_8_509));
   XNOR2_X1 i_8_383 (.A(n_8_509), .B(n_8_449), .ZN(n_8_510));
   OR2_X1 i_8_593 (.A1(n_8_509), .A2(n_58), .ZN(n_8_511));
   XNOR2_X1 i_8_386 (.A(n_8_509), .B(n_58), .ZN(n_8_512));
   NAND3_X1 i_8_394 (.A1(n_8_490), .A2(n_8_491), .A3(n_8_492), .ZN(n_8_513));
   NAND2_X1 i_8_375 (.A1(n_8_460), .A2(m[7]), .ZN(n_8_514));
   NAND2_X1 i_8_416 (.A1(n_8_411), .A2(n_8_415), .ZN(n_8_515));
   NAND2_X1 i_8_447 (.A1(n_8_413), .A2(n_8_414), .ZN(n_8_516));
   NAND2_X1 i_8_448 (.A1(n_8_460), .A2(m[7]), .ZN(n_8_517));
   NAND3_X1 i_8_604 (.A1(n_8_515), .A2(n_8_516), .A3(n_8_517), .ZN(n_8_518));
   NAND2_X1 i_8_250 (.A1(n_8_478), .A2(n_8_477), .ZN(n_8_519));
   INV_X1 i_8_258 (.A(n_8_519), .ZN(n_8_520));
   NAND2_X1 i_8_441 (.A1(n_8_438), .A2(n_8_433), .ZN(n_8_521));
   NAND2_X1 i_8_473 (.A1(n_8_450), .A2(n_8_434), .ZN(n_8_522));
   NAND3_X1 i_8_480 (.A1(n_8_521), .A2(n_8_522), .A3(n_8_424), .ZN(n_128));
   INV_X1 i_8_414 (.A(n_8_416), .ZN(n_8_523));
   NAND3_X1 i_8_442 (.A1(n_8_498), .A2(n_8_499), .A3(n_8_500), .ZN(n_8_524));
   INV_X1 i_8_496 (.A(n_60), .ZN(n_8_525));
   NAND2_X1 i_8_595 (.A1(n_8_500), .A2(n_8_525), .ZN(n_8_526));
   INV_X1 i_8_596 (.A(n_8_526), .ZN(n_8_527));
   NAND3_X1 i_8_597 (.A1(n_8_499), .A2(n_8_498), .A3(n_8_527), .ZN(n_8_528));
   INV_X1 i_8_401 (.A(n_8_528), .ZN(n_8_529));
   INV_X1 i_8_543 (.A(n_8_505), .ZN(n_8_530));
   NAND2_X1 i_8_489 (.A1(n_8_530), .A2(n_8_508), .ZN(n_8_531));
   XNOR2_X1 i_8_521 (.A(n_8_506), .B(n_8_507), .ZN(n_8_532));
   OAI21_X1 i_8_538 (.A(n_8_531), .B1(n_8_532), .B2(n_8_530), .ZN(n_8_533));
   NAND3_X1 i_8_472 (.A1(n_8_429), .A2(n_8_430), .A3(n_8_431), .ZN(n_129));
   INV_X1 i_8_598 (.A(m[7]), .ZN(n_8_534));
   NAND2_X1 i_8_607 (.A1(n_8_431), .A2(n_8_534), .ZN(n_8_535));
   INV_X1 i_8_608 (.A(n_8_535), .ZN(n_8_536));
   NAND3_X1 i_8_609 (.A1(n_8_429), .A2(n_8_430), .A3(n_8_536), .ZN(n_8_537));
   INV_X1 i_8_610 (.A(n_8_537), .ZN(n_8_538));
   NAND2_X1 i_8_481 (.A1(n_8_439), .A2(n_8_433), .ZN(n_8_539));
   NAND2_X1 i_8_483 (.A1(n_8_456), .A2(n_8_434), .ZN(n_8_540));
   NAND2_X1 i_8_603 (.A1(n_8_456), .A2(n_8_434), .ZN(n_8_541));
   NAND2_X1 i_8_611 (.A1(n_8_439), .A2(n_8_433), .ZN(n_8_542));
   NAND3_X1 i_8_612 (.A1(n_8_541), .A2(n_8_542), .A3(n_8_428), .ZN(n_8_543));
   NAND2_X1 i_8_560 (.A1(n_8_425), .A2(n_8_426), .ZN(n_8_544));
   NAND2_X1 i_8_570 (.A1(n_8_544), .A2(n_58), .ZN(n_8_545));
   NOR2_X1 i_8_573 (.A1(n_8_544), .A2(n_58), .ZN(n_8_546));
   NOR2_X1 i_8_574 (.A1(n_8_544), .A2(m[4]), .ZN(n_8_547));
   XNOR2_X1 i_8_576 (.A(n_130), .B(m[4]), .ZN(n_8_548));
   NAND2_X1 i_8_575 (.A1(n_8_425), .A2(n_8_426), .ZN(n_130));
   NAND3_X1 i_8_490 (.A1(n_8_501), .A2(n_8_502), .A3(n_8_503), .ZN(n_8_549));
   NAND2_X1 i_8_492 (.A1(n_8_553), .A2(n_55), .ZN(n_8_550));
   NAND2_X1 i_8_497 (.A1(n_8_549), .A2(m[9]), .ZN(n_8_551));
   NOR2_X1 i_8_498 (.A1(n_8_549), .A2(m[9]), .ZN(n_8_552));
   NAND3_X1 i_8_499 (.A1(n_8_501), .A2(n_8_502), .A3(n_8_503), .ZN(n_8_553));
   NAND2_X1 i_8_500 (.A1(n_8_452), .A2(n_8_434), .ZN(n_8_554));
   NAND2_X1 i_8_259 (.A1(n_8_443), .A2(n_8_444), .ZN(n_8_555));
   NAND2_X1 i_8_526 (.A1(n_8_443), .A2(n_8_444), .ZN(n_8_556));
   NAND2_X1 i_8_527 (.A1(n_8_452), .A2(n_8_434), .ZN(n_8_557));
   XNOR2_X1 i_8_581 (.A(n_8_454), .B(n_8_451), .ZN(n_8_558));
   NAND2_X1 i_8_582 (.A1(n_8_558), .A2(n_8_434), .ZN(n_8_559));
   NAND2_X1 i_8_475 (.A1(n_8_563), .A2(n_8_434), .ZN(n_8_560));
   NAND2_X1 i_8_479 (.A1(n_8_463), .A2(n_8_465), .ZN(n_8_561));
   NAND2_X1 i_8_617 (.A1(n_8_463), .A2(n_8_465), .ZN(n_8_562));
   NAND3_X1 i_8_618 (.A1(n_8_565), .A2(n_8_562), .A3(n_8_427), .ZN(n_131));
   XNOR2_X1 i_8_580 (.A(n_8_448), .B(n_8_453), .ZN(n_8_563));
   XNOR2_X1 i_8_606 (.A(n_8_448), .B(n_8_453), .ZN(n_8_564));
   NAND2_X1 i_8_619 (.A1(n_8_564), .A2(n_8_434), .ZN(n_8_565));
   NAND3_X1 i_8_614 (.A1(n_8_487), .A2(n_8_488), .A3(n_8_489), .ZN(n_8_566));
   XNOR2_X1 i_8_615 (.A(n_8_566), .B(m[3]), .ZN(n_8_567));
   NOR2_X1 i_8_616 (.A1(n_8_566), .A2(m[3]), .ZN(n_8_568));
   NAND3_X1 i_8_540 (.A1(n_8_487), .A2(n_8_488), .A3(n_8_489), .ZN(n_8_569));
   NAND3_X1 i_8_613 (.A1(n_8_556), .A2(n_8_557), .A3(n_8_432), .ZN(n_8_570));
   XNOR2_X1 i_8_620 (.A(n_8_570), .B(n_60), .ZN(n_8_571));
   NAND3_X1 i_8_621 (.A1(n_8_556), .A2(n_8_557), .A3(n_8_432), .ZN(n_132));
   INV_X1 i_8_53 (.A(m[6]), .ZN(n_8_572));
   XNOR2_X1 i_8_67 (.A(n_8_543), .B(n_8_572), .ZN(n_8_573));
   NAND2_X1 i_8_72 (.A1(n_8_469), .A2(n_8_421), .ZN(n_8_574));
   INV_X1 i_8_74 (.A(n_8_574), .ZN(n_8_575));
   AOI22_X1 i_8_82 (.A1(n_8_420), .A2(n_8_575), .B1(n_8_412), .B2(n_8_469), 
      .ZN(n_8_576));
   NAND2_X1 i_8_83 (.A1(n_8_573), .A2(n_8_576), .ZN(n_8_577));
   NAND2_X1 i_8_300 (.A1(n_8_460), .A2(n_69), .ZN(n_8_578));
   NAND3_X1 i_8_322 (.A1(n_8_429), .A2(n_8_430), .A3(n_8_445), .ZN(n_8_579));
   NAND2_X1 i_8_345 (.A1(n_8_578), .A2(n_8_579), .ZN(n_8_580));
   NAND3_X1 i_8_488 (.A1(n_8_539), .A2(n_8_540), .A3(n_8_428), .ZN(n_133));
   INV_X1 i_8_493 (.A(m[6]), .ZN(n_8_581));
   NAND2_X1 i_8_494 (.A1(n_8_428), .A2(n_8_581), .ZN(n_8_582));
   INV_X1 i_8_532 (.A(n_8_582), .ZN(n_8_583));
   NAND3_X1 i_8_587 (.A1(n_8_540), .A2(n_8_539), .A3(n_8_583), .ZN(n_8_584));
   INV_X1 i_8_589 (.A(n_8_584), .ZN(n_8_585));
   NAND3_X1 i_8_541 (.A1(n_8_495), .A2(n_8_496), .A3(n_8_497), .ZN(n_8_586));
   XNOR2_X1 i_8_542 (.A(n_8_586), .B(n_69), .ZN(n_8_587));
   NAND2_X1 i_8_544 (.A1(n_8_586), .A2(n_69), .ZN(n_8_588));
   XNOR2_X1 i_8_555 (.A(n_8_586), .B(m[7]), .ZN(n_8_589));
   OR2_X1 i_8_559 (.A1(n_8_586), .A2(m[7]), .ZN(n_8_590));
   NAND2_X1 i_8_594 (.A1(n_8_586), .A2(m[7]), .ZN(n_8_591));
   NAND3_X1 i_8_605 (.A1(n_8_495), .A2(n_8_496), .A3(n_8_497), .ZN(n_8_592));
endmodule

module Partial_Full_Adder__0_249(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_253(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_257(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_261(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_265(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_269(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_273(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_277(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_281(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_285(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   INV_X1 i_0_0 (.A(n_0_2), .ZN(G));
   INV_X1 i_0_6 (.A(A), .ZN(n_0_0));
   INV_X1 i_0_7 (.A(B), .ZN(n_0_1));
   NAND2_X1 i_0_2 (.A1(B), .A2(A), .ZN(n_0_2));
   AOI22_X1 i_0_3 (.A1(n_0_1), .A2(n_0_0), .B1(B), .B2(A), .ZN(P));
endmodule

module Partial_Full_Adder__0_289(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;
   wire n_0_1;

   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
   INV_X1 i_0_0 (.A(B), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(A), .ZN(n_0_1));
   OAI22_X1 i_0_4 (.A1(n_0_0), .A2(A), .B1(B), .B2(n_0_1), .ZN(P));
endmodule

module Partial_Full_Adder__0_293(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(P));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(A), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(B), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(B), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(A), .ZN(n_0_3));
   XOR2_X1 i_1_0 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_297(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   INV_X1 i_0_0 (.A(A), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(B), .B(n_0_0), .ZN(P));
   XOR2_X1 i_1_0 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_301(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   INV_X1 i_0_0 (.A(A), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(B), .B(n_0_0), .ZN(P));
   XOR2_X1 i_1_0 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_305(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;

   INV_X1 i_0_0 (.A(A), .ZN(n_0_0));
   OAI21_X1 i_0_1 (.A(n_0_1), .B1(B), .B2(n_0_2), .ZN(P));
   NAND2_X1 i_0_2 (.A1(B), .A2(n_0_0), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A), .ZN(n_0_2));
   NAND2_X1 i_1_0 (.A1(n_1_0), .A2(n_1_2), .ZN(S));
   NAND2_X1 i_1_1 (.A1(n_1_1), .A2(P), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(Cin), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(Cin), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(P), .ZN(n_1_3));
   AND2_X1 i_2_0 (.A1(B), .A2(A), .ZN(G));
endmodule

module Partial_Full_Adder(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XNOR2_X1 i_0_0 (.A(B), .B(A), .ZN(n_0_0));
   XNOR2_X1 i_0_1 (.A(Cin), .B(n_0_0), .ZN(S));
endmodule

module Carry_Look_Ahead(A, B, Cin, S);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]S;

   wire c1;
   wire c10;
   wire n_0_0;
   wire n_0_1;
   wire c11;
   wire n_1_0;
   wire n_1_1;
   wire c12;
   wire n_2_0;
   wire n_2_1;
   wire c13;
   wire n_3_0;
   wire n_3_1;
   wire n_6_0;
   wire c7;
   wire n_6_1;
   wire c6;
   wire n_6_2;
   wire c5;
   wire n_6_3;
   wire c4;
   wire n_6_4;
   wire c3;
   wire n_6_5;
   wire c2;
   wire n_6_6;
   wire c9;
   wire n_6_7;
   wire n_6_8;
   wire c8;
   wire c15;
   wire n_4_0;
   wire n_4_1;
   wire n_4_2;
   wire n_4_3;
   wire n_4_4;
   wire c14;
   wire n_5_0;
   wire n_5_1;

   Partial_Full_Adder__0_249 PFA1 (.A(A[0]), .B(B[0]), .Cin(), .S(S[0]), .P(), 
      .G(c1));
   Partial_Full_Adder__0_253 PFA2 (.A(A[1]), .B(B[1]), .Cin(c1), .S(S[1]), 
      .P(n_1), .G(n_0));
   Partial_Full_Adder__0_257 PFA3 (.A(A[2]), .B(B[2]), .Cin(c2), .S(S[2]), 
      .P(n_3), .G(n_2));
   Partial_Full_Adder__0_261 PFA4 (.A(A[3]), .B(B[3]), .Cin(c3), .S(S[3]), 
      .P(n_5), .G(n_4));
   Partial_Full_Adder__0_265 PFA5 (.A(A[4]), .B(B[4]), .Cin(c4), .S(S[4]), 
      .P(n_7), .G(n_6));
   Partial_Full_Adder__0_269 PFA6 (.A(A[5]), .B(B[5]), .Cin(c5), .S(S[5]), 
      .P(n_9), .G(n_8));
   Partial_Full_Adder__0_273 PFA7 (.A(A[6]), .B(B[6]), .Cin(c6), .S(S[6]), 
      .P(n_11), .G(n_10));
   Partial_Full_Adder__0_277 PFA8 (.A(A[7]), .B(B[7]), .Cin(c7), .S(S[7]), 
      .P(n_13), .G(n_12));
   Partial_Full_Adder__0_281 PFA9 (.A(A[8]), .B(B[8]), .Cin(c8), .S(S[8]), 
      .P(n_15), .G(n_14));
   Partial_Full_Adder__0_285 PFA10 (.A(A[9]), .B(B[9]), .Cin(c9), .S(S[9]), 
      .P(n_17), .G(n_16));
   Partial_Full_Adder__0_289 PFA11 (.A(A[10]), .B(B[10]), .Cin(c10), .S(S[10]), 
      .P(n_19), .G(n_18));
   Partial_Full_Adder__0_293 PFA12 (.A(A[11]), .B(B[11]), .Cin(c11), .S(S[11]), 
      .P(n_21), .G(n_20));
   Partial_Full_Adder__0_297 PFA13 (.A(A[12]), .B(B[12]), .Cin(c12), .S(S[12]), 
      .P(n_23), .G(n_22));
   Partial_Full_Adder__0_301 PFA14 (.A(A[13]), .B(B[13]), .Cin(c13), .S(S[13]), 
      .P(n_25), .G(n_24));
   Partial_Full_Adder__0_305 PFA15 (.A(A[14]), .B(B[14]), .Cin(c14), .S(S[14]), 
      .P(n_27), .G(n_26));
   Partial_Full_Adder PFA16 (.A(A[15]), .B(B[15]), .Cin(c15), .S(S[15]), .P(), 
      .G());
   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_1), .ZN(c10));
   NAND2_X1 i_0_1 (.A1(n_17), .A2(c9), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_16), .ZN(n_0_1));
   NAND2_X1 i_1_0 (.A1(n_1_0), .A2(n_1_1), .ZN(c11));
   NAND2_X1 i_1_1 (.A1(c10), .A2(n_19), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_18), .ZN(n_1_1));
   NAND2_X1 i_2_0 (.A1(n_2_0), .A2(n_2_1), .ZN(c12));
   NAND2_X1 i_2_1 (.A1(n_21), .A2(c11), .ZN(n_2_0));
   INV_X1 i_2_2 (.A(n_20), .ZN(n_2_1));
   NAND2_X1 i_3_0 (.A1(n_3_0), .A2(n_3_1), .ZN(c13));
   NAND2_X1 i_3_1 (.A1(c12), .A2(n_23), .ZN(n_3_0));
   INV_X1 i_3_2 (.A(n_22), .ZN(n_3_1));
   AOI21_X1 i_6_0 (.A(n_12), .B1(n_13), .B2(c7), .ZN(n_6_0));
   INV_X1 i_6_1 (.A(n_6_1), .ZN(c7));
   AOI21_X1 i_6_2 (.A(n_10), .B1(n_11), .B2(c6), .ZN(n_6_1));
   INV_X1 i_6_3 (.A(n_6_2), .ZN(c6));
   AOI21_X1 i_6_4 (.A(n_8), .B1(n_9), .B2(c5), .ZN(n_6_2));
   INV_X1 i_6_5 (.A(n_6_3), .ZN(c5));
   AOI21_X1 i_6_6 (.A(n_6), .B1(n_7), .B2(c4), .ZN(n_6_3));
   INV_X1 i_6_7 (.A(n_6_4), .ZN(c4));
   AOI21_X1 i_6_8 (.A(n_4), .B1(n_5), .B2(c3), .ZN(n_6_4));
   INV_X1 i_6_9 (.A(n_6_5), .ZN(c3));
   AOI21_X1 i_6_10 (.A(n_2), .B1(n_3), .B2(c2), .ZN(n_6_5));
   INV_X1 i_6_11 (.A(n_6_6), .ZN(c2));
   AOI21_X1 i_6_12 (.A(n_0), .B1(c1), .B2(n_1), .ZN(n_6_6));
   NAND2_X1 i_6_13 (.A1(n_6_7), .A2(n_6_8), .ZN(c9));
   NAND2_X1 i_6_14 (.A1(n_15), .A2(c8), .ZN(n_6_7));
   INV_X1 i_6_15 (.A(n_14), .ZN(n_6_8));
   INV_X1 i_6_16 (.A(n_6_0), .ZN(c8));
   NAND2_X1 i_4_0 (.A1(n_4_0), .A2(n_4_4), .ZN(c15));
   NAND2_X1 i_4_1 (.A1(n_4_1), .A2(n_27), .ZN(n_4_0));
   NAND2_X1 i_4_2 (.A1(n_4_2), .A2(n_4_3), .ZN(n_4_1));
   NAND2_X1 i_4_3 (.A1(n_25), .A2(c13), .ZN(n_4_2));
   INV_X1 i_4_4 (.A(n_24), .ZN(n_4_3));
   INV_X1 i_4_5 (.A(n_26), .ZN(n_4_4));
   NAND2_X1 i_5_0 (.A1(n_5_0), .A2(n_5_1), .ZN(c14));
   NAND2_X1 i_5_1 (.A1(n_25), .A2(c13), .ZN(n_5_0));
   INV_X1 i_5_2 (.A(n_24), .ZN(n_5_1));
endmodule

module Interpolation_Logic(Un, Uz, DivResult, EN, Uk);
   input [15:0]Un;
   input [15:0]Uz;
   input [15:0]DivResult;
   input EN;
   output [15:0]Uk;

   wire [15:0]UnComp;
   wire [15:0]Uz_Un;
   wire [15:0]secondOperand;
   wire [15:0]temp;

   Carry_Look_Ahead__0_710 add1 (.A(temp), .B(), .Cin(), .S({UnComp[15], 
      UnComp[14], UnComp[13], UnComp[12], UnComp[11], UnComp[10], UnComp[9], 
      UnComp[8], UnComp[7], UnComp[6], UnComp[5], UnComp[4], UnComp[3], 
      UnComp[2], UnComp[1], uc_0}));
   Carry_Look_Ahead__0_791 Sub (.A(Uz), .B({UnComp[15], UnComp[14], UnComp[13], 
      UnComp[12], UnComp[11], UnComp[10], UnComp[9], UnComp[8], UnComp[7], 
      UnComp[6], UnComp[5], UnComp[4], UnComp[3], UnComp[2], UnComp[1], Un[0]}), 
      .Cin(), .S(Uz_Un));
   booth_multiplier mul (.m(DivResult), .r(Uz_Un), .result(secondOperand), 
      .overflow());
   Carry_Look_Ahead add (.A(Un), .B(secondOperand), .Cin(), .S(Uk));
   INV_X1 i_0_0 (.A(Un[0]), .ZN(temp[0]));
   INV_X1 i_0_1 (.A(Un[1]), .ZN(temp[1]));
   INV_X1 i_0_2 (.A(Un[2]), .ZN(temp[2]));
   INV_X1 i_0_3 (.A(Un[3]), .ZN(temp[3]));
   INV_X1 i_0_4 (.A(Un[4]), .ZN(temp[4]));
   INV_X1 i_0_5 (.A(Un[5]), .ZN(temp[5]));
   INV_X1 i_0_6 (.A(Un[6]), .ZN(temp[6]));
   INV_X1 i_0_7 (.A(Un[7]), .ZN(temp[7]));
   INV_X1 i_0_8 (.A(Un[8]), .ZN(temp[8]));
   INV_X1 i_0_9 (.A(Un[9]), .ZN(temp[9]));
   INV_X1 i_0_10 (.A(Un[10]), .ZN(temp[10]));
   INV_X1 i_0_11 (.A(Un[11]), .ZN(temp[11]));
   INV_X1 i_0_12 (.A(Un[12]), .ZN(temp[12]));
   INV_X1 i_0_13 (.A(Un[13]), .ZN(temp[13]));
   INV_X1 i_0_14 (.A(Un[14]), .ZN(temp[14]));
   INV_X1 i_0_15 (.A(Un[15]), .ZN(temp[15]));
endmodule

module Interpolation(Tk, Uz, Un, Tz, CLK, reset, DivFlag, shiftFlag, DivDoneFlag, 
      Uk);
   input [15:0]Tk;
   input [15:0]Uz;
   input [15:0]Un;
   input [15:0]Tz;
   input CLK;
   input reset;
   input DivFlag;
   input shiftFlag;
   output DivDoneFlag;
   output [15:0]Uk;

   wire [15:0]Div_Output;
   wire [15:0]Tz_RegTemp;
   wire [15:0]Tn_RegTemp;
   wire [15:0]Div_Output_Reg;
   wire [15:0]Tn_Reg;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;

   Interpolation_Devision Dk (.Tk(Tk), .Tz(Tz), .Tn(Tn_Reg), .CLK(CLK), .reset(
      reset), .EN(DivFlag), .Done(DivDoneFlag), .DivOut(Div_Output));
   reg__0_811 Reg_Tz (.D(Tz), .load(), .Clk(CLK), .Q(Tz_RegTemp), .rst(reset));
   reg__0_831 Reg_Tn (.D(Tz_RegTemp), .load(shiftFlag), .Clk(CLK), .Q(Tn_RegTemp), 
      .rst(reset));
   \reg  DivOut_Reg (.D(Div_Output), .load(DivDoneFlag), .Clk(CLK), .Q(
      Div_Output_Reg), .rst(reset));
   Interpolation_Logic L1 (.Un(Un), .Uz(Uz), .DivResult(Div_Output_Reg), .EN(), 
      .Uk(Uk));
   DLH_X1 \Tn_Reg_reg[15]  (.D(n_0_15), .G(n_0_16), .Q(Tn_Reg[15]));
   DLH_X1 \Tn_Reg_reg[14]  (.D(n_0_14), .G(n_0_16), .Q(Tn_Reg[14]));
   DLH_X1 \Tn_Reg_reg[13]  (.D(n_0_13), .G(n_0_16), .Q(Tn_Reg[13]));
   DLH_X1 \Tn_Reg_reg[12]  (.D(n_0_12), .G(n_0_16), .Q(Tn_Reg[12]));
   DLH_X1 \Tn_Reg_reg[11]  (.D(n_0_11), .G(n_0_16), .Q(Tn_Reg[11]));
   DLH_X1 \Tn_Reg_reg[10]  (.D(n_0_10), .G(n_0_16), .Q(Tn_Reg[10]));
   DLH_X1 \Tn_Reg_reg[9]  (.D(n_0_9), .G(n_0_16), .Q(Tn_Reg[9]));
   DLH_X1 \Tn_Reg_reg[8]  (.D(n_0_8), .G(n_0_16), .Q(Tn_Reg[8]));
   DLH_X1 \Tn_Reg_reg[7]  (.D(n_0_7), .G(n_0_16), .Q(Tn_Reg[7]));
   DLH_X1 \Tn_Reg_reg[6]  (.D(n_0_6), .G(n_0_16), .Q(Tn_Reg[6]));
   DLH_X1 \Tn_Reg_reg[5]  (.D(n_0_5), .G(n_0_16), .Q(Tn_Reg[5]));
   DLH_X1 \Tn_Reg_reg[4]  (.D(n_0_4), .G(n_0_16), .Q(Tn_Reg[4]));
   DLH_X1 \Tn_Reg_reg[3]  (.D(n_0_3), .G(n_0_16), .Q(Tn_Reg[3]));
   DLH_X1 \Tn_Reg_reg[2]  (.D(n_0_2), .G(n_0_16), .Q(Tn_Reg[2]));
   DLH_X1 \Tn_Reg_reg[1]  (.D(n_0_1), .G(n_0_16), .Q(Tn_Reg[1]));
   DLH_X1 \Tn_Reg_reg[0]  (.D(n_0_0), .G(n_0_16), .Q(Tn_Reg[0]));
   AND2_X1 i_0_0_0 (.A1(shiftFlag), .A2(Tn_RegTemp[0]), .ZN(n_0_0));
   AND2_X1 i_0_0_1 (.A1(Tn_RegTemp[1]), .A2(shiftFlag), .ZN(n_0_1));
   AND2_X1 i_0_0_2 (.A1(Tn_RegTemp[2]), .A2(shiftFlag), .ZN(n_0_2));
   AND2_X1 i_0_0_3 (.A1(Tn_RegTemp[3]), .A2(shiftFlag), .ZN(n_0_3));
   AND2_X1 i_0_0_4 (.A1(Tn_RegTemp[4]), .A2(shiftFlag), .ZN(n_0_4));
   AND2_X1 i_0_0_5 (.A1(Tn_RegTemp[5]), .A2(shiftFlag), .ZN(n_0_5));
   AND2_X1 i_0_0_6 (.A1(Tn_RegTemp[6]), .A2(shiftFlag), .ZN(n_0_6));
   AND2_X1 i_0_0_7 (.A1(Tn_RegTemp[7]), .A2(shiftFlag), .ZN(n_0_7));
   AND2_X1 i_0_0_8 (.A1(Tn_RegTemp[8]), .A2(shiftFlag), .ZN(n_0_8));
   AND2_X1 i_0_0_9 (.A1(Tn_RegTemp[9]), .A2(shiftFlag), .ZN(n_0_9));
   AND2_X1 i_0_0_10 (.A1(Tn_RegTemp[10]), .A2(shiftFlag), .ZN(n_0_10));
   AND2_X1 i_0_0_11 (.A1(Tn_RegTemp[11]), .A2(shiftFlag), .ZN(n_0_11));
   AND2_X1 i_0_0_12 (.A1(Tn_RegTemp[12]), .A2(shiftFlag), .ZN(n_0_12));
   AND2_X1 i_0_0_13 (.A1(Tn_RegTemp[13]), .A2(shiftFlag), .ZN(n_0_13));
   AND2_X1 i_0_0_14 (.A1(Tn_RegTemp[14]), .A2(shiftFlag), .ZN(n_0_14));
   AND2_X1 i_0_0_15 (.A1(Tn_RegTemp[15]), .A2(shiftFlag), .ZN(n_0_15));
   OR2_X1 i_0_0_16 (.A1(reset), .A2(shiftFlag), .ZN(n_0_16));
endmodule
