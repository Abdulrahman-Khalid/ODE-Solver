/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 07:15:46 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2853951044 */

module FullAdder__1_476(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__1_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_347(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_344(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(in1), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_341(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__1_477(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__1_476 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__1_383 muxx_1_muxx_j (.sel(A[0]), .in1(A[1]), .in2(), .i1(), .i2(), 
      .out1(sum[1]), .Carry(n_5));
   mux__1_380 muxx_2_muxx_j (.sel(n_5), .in1(A[2]), .in2(), .i1(), .i2(), 
      .out1(sum[2]), .Carry(n_9));
   mux__1_377 muxx_3_muxx_j (.sel(n_9), .in1(A[3]), .in2(), .i1(), .i2(), 
      .out1(sum[3]), .Carry(n_0));
   mux__1_374 muxx_4_muxx_j (.sel(n_0), .in1(A[4]), .in2(), .i1(), .i2(), 
      .out1(sum[4]), .Carry(n_1));
   mux__1_371 muxx_5_muxx_j (.sel(n_1), .in1(A[5]), .in2(), .i1(), .i2(), 
      .out1(sum[5]), .Carry(n_2));
   mux__1_368 muxx_6_muxx_j (.sel(n_2), .in1(A[6]), .in2(), .i1(), .i2(), 
      .out1(sum[6]), .Carry(n_3));
   mux__1_365 muxx_7_muxx_j (.sel(n_3), .in1(A[7]), .in2(), .i1(), .i2(), 
      .out1(sum[7]), .Carry(n_4));
   mux__1_362 muxx_8_muxx_j (.sel(n_4), .in1(A[8]), .in2(), .i1(), .i2(), 
      .out1(sum[8]), .Carry(n_6));
   mux__1_359 muxx_9_muxx_j (.sel(n_6), .in1(A[9]), .in2(), .i1(), .i2(), 
      .out1(sum[9]), .Carry(n_7));
   mux__1_356 muxx_10_muxx_j (.sel(n_7), .in1(A[10]), .in2(), .i1(), .i2(), 
      .out1(sum[10]), .Carry(n_8));
   mux__1_353 muxx_11_muxx_j (.sel(n_8), .in1(A[11]), .in2(), .i1(), .i2(), 
      .out1(sum[11]), .Carry(n_10));
   mux__1_350 muxx_12_muxx_j (.sel(n_10), .in1(A[12]), .in2(), .i1(), .i2(), 
      .out1(sum[12]), .Carry(n_11));
   mux__1_347 muxx_13_muxx_j (.sel(n_11), .in1(A[13]), .in2(), .i1(), .i2(), 
      .out1(sum[13]), .Carry(n_12));
   mux__1_344 muxx_14_muxx_j (.sel(n_12), .in1(A[14]), .in2(), .i1(), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__1_341 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__1_327(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__1_321(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__1_315(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__1_312(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_309(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_306(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_303(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_300(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_297(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_294(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_291(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_288(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_285(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__1_282(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__1_219(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__1_216(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__1_213(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__1_210(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__1_207(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__1_204(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_201(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__1_198(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__1_334(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__1_327 FA_15_FA0_i (.in1(), .in2(B[15]), .Ci(), .S(n_2), .Co());
   FullAdder__1_321 FA_14_FA0_i (.in1(), .in2(B[14]), .Ci(), .S(n_6), .Co());
   FullAdder__1_315 FA_13_FA0_i (.in1(), .in2(B[13]), .Ci(), .S(n_10), .Co());
   FullAdder__1_312 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__1_309 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__1_306 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__1_303 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__1_300 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__1_297 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__1_294 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__1_291 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__1_288 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__1_285 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_0), .Co(n_29));
   FullAdder__1_282 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_1));
   mux__1_219 muxx_8_muxx_j (.sel(n_1), .in1(n_0), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_3));
   mux__1_216 muxx_9_muxx_j (.sel(n_3), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_4));
   mux__1_213 muxx_10_muxx_j (.sel(n_4), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_5));
   mux__1_210 muxx_11_muxx_j (.sel(n_5), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_7));
   mux__1_207 muxx_12_muxx_j (.sel(n_7), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_8));
   mux__1_204 muxx_13_muxx_j (.sel(n_8), .in1(n_10), .in2(), .i1(B[13]), .i2(), 
      .out1(sum[13]), .Carry(n_9));
   mux__1_201 muxx_14_muxx_j (.sel(n_9), .in1(n_6), .in2(), .i1(B[14]), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__1_198 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__1_334 u1 (.A({uc_0, uc_1, uc_2, notplus[12], notplus[11], 
      notplus[10], notplus[9], notplus[8], notplus[7], uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9}), .B({firstVal[15], firstVal[14], firstVal[13], 
      firstVal[12], firstVal[11], firstVal[10], firstVal[9], firstVal[8], 
      firstVal[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16}), .Cin(), 
      .sum({n_0, sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
      sum[7], uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23}), .overFlow());
   NOR4_X1 i_0_0 (.A1(firstVal[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), 
      .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(firstVal[6]), .A4(firstVal[5]), 
      .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(firstVal[4]), .A2(firstVal[3]), .A3(firstVal[2]), .A4(
      firstVal[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
endmodule

module counterMux(counter, resetdata, dataIn, start, load, reset, universalReset, 
      continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(counter[0]), .A2(n_0_0), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(counter[1]), .A2(n_0_0), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(counter[2]), .A2(n_0_0), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(counter[3]), .A2(n_0_0), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(counter[4]), .A2(n_0_0), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(counter[5]), .A2(n_0_0), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(counter[6]), .A2(n_0_0), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(counter[7]), .A2(n_0_0), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(counter[8]), .A2(n_0_0), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(counter[9]), .A2(n_0_0), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(counter[10]), .A2(n_0_0), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(counter[11]), .A2(n_0_0), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(counter[12]), .A2(n_0_0), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(counter[13]), .A2(n_0_0), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(counter[14]), .A2(n_0_0), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(counter[15]), .A2(n_0_0), .ZN(result[15]));
   NOR2_X1 i_0_16 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
endmodule

module reg__1_59(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]muxOut;
   wire activate;

   Addition1__1_477 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   comparator compare (.firstVal(dataOut), .secondVal({uc_0, uc_1, uc_2, 
      offset[12], offset[11], offset[10], offset[9], offset[8], offset[7], uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .done(done), .firstBigger(), 
      .firstSmaller());
   counterMux muxing (.counter(incremented), .resetdata(), .dataIn(), .start(), 
      .load(), .reset(done), .universalReset(universalReset), .continue(), 
      .result(muxOut));
   reg__1_59 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   OR3_X1 i_0_0 (.A1(universalReset), .A2(done), .A3(enable), .ZN(activate));
endmodule

module FullAdder__14_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__14_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__14_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__14_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__14_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__14_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__14_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__14_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__14_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__14_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__14_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__14_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__14_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__14_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__14_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__14_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__14_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__14_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__14_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__14_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__14_308(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_305(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_302(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_299(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_296(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_293(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_290(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_287(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_284(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_281(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_275(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__14_215(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_212(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_209(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_206(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_203(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_200(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_0_0 (.A(in1), .B(sel), .Z(out1));
   AND2_X1 i_0_1 (.A1(sel), .A2(in1), .ZN(Carry));
endmodule

module mux__14_197(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_0_0 (.A(in1), .B(sel), .Z(out1));
   AND2_X1 i_0_1 (.A1(sel), .A2(in1), .ZN(Carry));
endmodule

module mux__14_194(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__14_328(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__14_308 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__14_305 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__14_302 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__14_299 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__14_296 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__14_293 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__14_290 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__14_287 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__14_284 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_1), 
      .Co(n_0));
   FullAdder__14_281 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_3), 
      .Co(n_2));
   FullAdder__14_275 FA_7_FA0_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_4));
   mux__14_215 muxx_8_muxx_j (.sel(n_4), .in1(n_3), .in2(n_1), .i1(n_2), 
      .i2(n_0), .out1(sum[8]), .Carry(n_5));
   mux__14_212 muxx_9_muxx_j (.sel(n_5), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_6));
   mux__14_209 muxx_10_muxx_j (.sel(n_6), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_7));
   mux__14_206 muxx_11_muxx_j (.sel(n_7), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_8));
   mux__14_203 muxx_12_muxx_j (.sel(n_8), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_9));
   mux__14_200 muxx_13_muxx_j (.sel(n_9), .in1(A[13]), .in2(), .i1(), .i2(), 
      .out1(sum[13]), .Carry(n_10));
   mux__14_197 muxx_14_muxx_j (.sel(n_10), .in1(A[14]), .in2(), .i1(), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__14_194 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__14_190(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_187(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_1 (.A(in1), .B(in2), .ZN(S));
endmodule

module FullAdder__14_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in2), .B(in1), .Z(S));
endmodule

module FullAdder__14_183(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_177(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_138(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_135(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_132(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_129(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_126(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_123(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_120(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_117(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_114(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_111(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_108(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_105(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__14_102(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__14_99(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_96(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_93(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_90(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_87(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_84(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_81(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__14_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_1_0 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module Addition1__14_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire S;
   wire Carry;

   FullAdder__14_190 FA0 (.in1(A[0]), .in2(B[0]), .Ci(), .S(sum[0]), .Co(n_0));
   FullAdder__14_187 FA_15_FA1_i (.in1(A[15]), .in2(B[15]), .Ci(), .S(S), .Co());
   FullAdder__14_185 FA_15_FA0_i (.in1(A[15]), .in2(B[15]), .Ci(), .S(n_2), 
      .Co());
   FullAdder__14_183 FA_14_FA1_i (.in1(A[14]), .in2(B[14]), .Ci(), .S(n_4), 
      .Co(n_3));
   FullAdder__14_180 FA_14_FA0_i (.in1(A[14]), .in2(B[14]), .Ci(), .S(n_6), 
      .Co(n_5));
   FullAdder__14_177 FA_13_FA1_i (.in1(A[13]), .in2(B[13]), .Ci(), .S(n_8), 
      .Co(n_7));
   FullAdder__14_174 FA_13_FA0_i (.in1(A[13]), .in2(B[13]), .Ci(), .S(n_10), 
      .Co(n_9));
   FullAdder__14_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__14_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__14_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__14_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__14_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__14_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__14_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__14_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__14_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__14_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_30), 
      .Co(n_29));
   FullAdder__14_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(n_32), 
      .Co(n_31));
   FullAdder__14_138 FA_7_FA0_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(n_34), 
      .Co(n_33));
   FullAdder__14_135 FA_6_FA1_i (.in1(A[6]), .in2(B[6]), .Ci(), .S(n_36), 
      .Co(n_35));
   FullAdder__14_132 FA_6_FA0_i (.in1(A[6]), .in2(B[6]), .Ci(), .S(n_38), 
      .Co(n_37));
   FullAdder__14_129 FA_5_FA1_i (.in1(A[5]), .in2(B[5]), .Ci(), .S(n_40), 
      .Co(n_39));
   FullAdder__14_126 FA_5_FA0_i (.in1(A[5]), .in2(B[5]), .Ci(), .S(n_42), 
      .Co(n_41));
   FullAdder__14_123 FA_4_FA1_i (.in1(A[4]), .in2(B[4]), .Ci(), .S(n_44), 
      .Co(n_43));
   FullAdder__14_120 FA_4_FA0_i (.in1(A[4]), .in2(B[4]), .Ci(), .S(n_46), 
      .Co(n_45));
   FullAdder__14_117 FA_3_FA1_i (.in1(A[3]), .in2(B[3]), .Ci(), .S(n_48), 
      .Co(n_47));
   FullAdder__14_114 FA_3_FA0_i (.in1(A[3]), .in2(B[3]), .Ci(), .S(n_50), 
      .Co(n_49));
   FullAdder__14_111 FA_2_FA1_i (.in1(A[2]), .in2(B[2]), .Ci(), .S(n_52), 
      .Co(n_51));
   FullAdder__14_108 FA_2_FA0_i (.in1(A[2]), .in2(B[2]), .Ci(), .S(n_54), 
      .Co(n_53));
   FullAdder__14_105 FA_1_FA1_i (.in1(A[1]), .in2(B[1]), .Ci(), .S(n_56), 
      .Co(n_55));
   FullAdder__14_102 FA_1_FA0_i (.in1(A[1]), .in2(B[1]), .Ci(), .S(n_58), 
      .Co(n_57));
   mux__14_99 muxx_1_muxx_j (.sel(n_0), .in1(n_58), .in2(n_56), .i1(n_57), 
      .i2(n_55), .out1(sum[1]), .Carry(n_59));
   mux__14_96 muxx_2_muxx_j (.sel(n_59), .in1(n_54), .in2(n_52), .i1(n_53), 
      .i2(n_51), .out1(sum[2]), .Carry(n_60));
   mux__14_93 muxx_3_muxx_j (.sel(n_60), .in1(n_50), .in2(n_48), .i1(n_49), 
      .i2(n_47), .out1(sum[3]), .Carry(n_61));
   mux__14_90 muxx_4_muxx_j (.sel(n_61), .in1(n_46), .in2(n_44), .i1(n_45), 
      .i2(n_43), .out1(sum[4]), .Carry(n_62));
   mux__14_87 muxx_5_muxx_j (.sel(n_62), .in1(n_42), .in2(n_40), .i1(n_41), 
      .i2(n_39), .out1(sum[5]), .Carry(n_63));
   mux__14_84 muxx_6_muxx_j (.sel(n_63), .in1(n_38), .in2(n_36), .i1(n_37), 
      .i2(n_35), .out1(sum[6]), .Carry(n_64));
   mux__14_81 muxx_7_muxx_j (.sel(n_64), .in1(n_34), .in2(n_32), .i1(n_33), 
      .i2(n_31), .out1(sum[7]), .Carry(n_65));
   mux__14_78 muxx_8_muxx_j (.sel(n_65), .in1(n_30), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_66));
   mux__14_75 muxx_9_muxx_j (.sel(n_66), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_67));
   mux__14_72 muxx_10_muxx_j (.sel(n_67), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_68));
   mux__14_69 muxx_11_muxx_j (.sel(n_68), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_69));
   mux__14_66 muxx_12_muxx_j (.sel(n_69), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_70));
   mux__14_63 muxx_13_muxx_j (.sel(n_70), .in1(n_10), .in2(n_8), .i1(n_9), 
      .i2(n_7), .out1(sum[13]), .Carry(n_1));
   mux__14_60 muxx_14_muxx_j (.sel(n_1), .in1(n_6), .in2(n_4), .i1(n_5), 
      .i2(n_3), .out1(sum[14]), .Carry(Carry));
   mux__14_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(S), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__14_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__14_191 u1 (.A(notplus), .B(firstVal), .Cin(), .sum({n_0, sum[14], 
      sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], sum[7], sum[6], sum[5], 
      sum[4], sum[3], sum[2], sum[1], sum[0]}), .overFlow());
   NOR4_X1 i_0_0 (.A1(sum[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(sum[6]), .A4(sum[5]), .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(sum[4]), .A2(sum[3]), .A3(sum[2]), .A4(sum[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_0 (.A(secondVal[0]), .ZN(notplus[0]));
   INV_X1 i_1_1 (.A(secondVal[1]), .ZN(notplus[1]));
   INV_X1 i_1_2 (.A(secondVal[2]), .ZN(notplus[2]));
   INV_X1 i_1_3 (.A(secondVal[3]), .ZN(notplus[3]));
   INV_X1 i_1_4 (.A(secondVal[4]), .ZN(notplus[4]));
   INV_X1 i_1_5 (.A(secondVal[5]), .ZN(notplus[5]));
   INV_X1 i_1_6 (.A(secondVal[6]), .ZN(notplus[6]));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
   INV_X1 i_1_13 (.A(secondVal[13]), .ZN(notplus[13]));
   INV_X1 i_1_14 (.A(secondVal[14]), .ZN(notplus[14]));
   INV_X1 i_1_15 (.A(secondVal[15]), .ZN(notplus[15]));
endmodule

module smallMux__14_53(loadAddress, CurrentCount, start, universalReset, 
      innerDone, continue, load, address);
   input [15:0]loadAddress;
   input [15:0]CurrentCount;
   input [15:0]start;
   input universalReset;
   input innerDone;
   input continue;
   input load;
   output [15:0]address;

   wire n_0_0;
   wire n_0_1;

   AND2_X1 i_0_0 (.A1(CurrentCount[0]), .A2(n_0_0), .ZN(address[0]));
   AND2_X1 i_0_1 (.A1(CurrentCount[1]), .A2(n_0_0), .ZN(address[1]));
   AND2_X1 i_0_2 (.A1(CurrentCount[2]), .A2(n_0_0), .ZN(address[2]));
   AND2_X1 i_0_3 (.A1(CurrentCount[3]), .A2(n_0_0), .ZN(address[3]));
   AND2_X1 i_0_4 (.A1(CurrentCount[4]), .A2(n_0_0), .ZN(address[4]));
   AND2_X1 i_0_5 (.A1(CurrentCount[5]), .A2(n_0_0), .ZN(address[5]));
   AND2_X1 i_0_6 (.A1(CurrentCount[6]), .A2(n_0_0), .ZN(address[6]));
   AND2_X1 i_0_7 (.A1(CurrentCount[7]), .A2(n_0_0), .ZN(address[7]));
   AND2_X1 i_0_8 (.A1(CurrentCount[8]), .A2(n_0_0), .ZN(address[8]));
   AND2_X1 i_0_9 (.A1(CurrentCount[9]), .A2(n_0_0), .ZN(address[9]));
   AND2_X1 i_0_10 (.A1(CurrentCount[10]), .A2(n_0_0), .ZN(address[10]));
   AND2_X1 i_0_11 (.A1(CurrentCount[11]), .A2(n_0_0), .ZN(address[11]));
   AND2_X1 i_0_12 (.A1(CurrentCount[12]), .A2(n_0_0), .ZN(address[12]));
   AND2_X1 i_0_13 (.A1(CurrentCount[13]), .A2(n_0_0), .ZN(address[13]));
   AND2_X1 i_0_14 (.A1(CurrentCount[14]), .A2(n_0_0), .ZN(address[14]));
   AND2_X1 i_0_15 (.A1(CurrentCount[15]), .A2(n_0_0), .ZN(address[15]));
   NOR2_X1 i_0_16 (.A1(n_0_1), .A2(universalReset), .ZN(n_0_0));
   NAND2_X1 i_0_17 (.A1(continue), .A2(innerDone), .ZN(n_0_1));
endmodule

module reg__14_49(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counterMux__14_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(n_0_0), .A2(counter[0]), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(counter[1]), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(counter[2]), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(counter[3]), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(counter[4]), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(counter[5]), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(counter[6]), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(counter[7]), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(counter[8]), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(counter[9]), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(counter[10]), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(counter[11]), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(counter[12]), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(counter[13]), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(counter[14]), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(counter[15]), .ZN(result[15]));
   INV_X1 i_0_16 (.A(universalReset), .ZN(n_0_0));
endmodule

module reg__14_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__1_478(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]plus;
   wire [15:0]newStart;
   wire [15:0]init;
   wire [15:0]muxOut;
   wire setNewstart;
   wire n_0_0;
   wire activate;
   wire n_0_1;
   wire n_0_2;

   Addition1__14_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   Addition1__14_328 u0 (.A({init[15], init[14], init[13], init[12], init[11], 
      init[10], init[9], init[8], init[7], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, 
      uc_6}), .B({uc_7, uc_8, uc_9, offset[12], offset[11], offset[10], 
      offset[9], offset[8], offset[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16}), .Cin(), .sum({plus[15], plus[14], plus[13], plus[12], plus[11], 
      plus[10], plus[9], plus[8], plus[7], uc_17, uc_18, uc_19, uc_20, uc_21, 
      uc_22, uc_23}), .overFlow());
   comparator__14_192 compare (.firstVal(dataOut), .secondVal({plus[15], 
      plus[14], plus[13], plus[12], plus[11], plus[10], plus[9], plus[8], 
      plus[7], init[6], init[5], init[4], init[3], init[2], init[1], init[0]}), 
      .done(done), .firstBigger(), .firstSmaller());
   smallMux__14_53 smallMux (.loadAddress(), .CurrentCount(dataOut), .start(), 
      .universalReset(universalReset), .innerDone(done), .continue(continue), 
      .load(), .address(newStart));
   reg__14_49 initialAdress (.D(newStart), .load(setNewstart), .Clk(CLK), 
      .Q(init), .rst(universalReset));
   counterMux__14_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(), .universalReset(universalReset), .continue(), 
      .result(muxOut));
   reg__14_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   INV_X1 i_0_0 (.A(n_0_0), .ZN(setNewstart));
   AOI21_X1 i_0_1 (.A(universalReset), .B1(done), .B2(continue), .ZN(n_0_0));
   OAI21_X1 i_0_2 (.A(n_0_2), .B1(n_0_1), .B2(done), .ZN(activate));
   INV_X1 i_0_3 (.A(enable), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(universalReset), .ZN(n_0_2));
endmodule

module FullAdder__15_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__15_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__15_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__15_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__15_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__15_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__15_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__15_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__15_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__15_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__15_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__15_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__15_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__15_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__15_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__15_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__15_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__15_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__15_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__15_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__15_308(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_305(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_302(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_299(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_296(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_293(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_290(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_287(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_284(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_281(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_275(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__15_215(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_212(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_209(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_206(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_203(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_200(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_0_0 (.A(in1), .B(sel), .Z(out1));
   AND2_X1 i_0_1 (.A1(sel), .A2(in1), .ZN(Carry));
endmodule

module mux__15_197(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_0_0 (.A(in1), .B(sel), .Z(out1));
   AND2_X1 i_0_1 (.A1(sel), .A2(in1), .ZN(Carry));
endmodule

module mux__15_194(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__15_328(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__15_308 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__15_305 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__15_302 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__15_299 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__15_296 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__15_293 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__15_290 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__15_287 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__15_284 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_1), 
      .Co(n_0));
   FullAdder__15_281 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_3), 
      .Co(n_2));
   FullAdder__15_275 FA_7_FA0_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_4));
   mux__15_215 muxx_8_muxx_j (.sel(n_4), .in1(n_3), .in2(n_1), .i1(n_2), 
      .i2(n_0), .out1(sum[8]), .Carry(n_5));
   mux__15_212 muxx_9_muxx_j (.sel(n_5), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_6));
   mux__15_209 muxx_10_muxx_j (.sel(n_6), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_7));
   mux__15_206 muxx_11_muxx_j (.sel(n_7), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_8));
   mux__15_203 muxx_12_muxx_j (.sel(n_8), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_9));
   mux__15_200 muxx_13_muxx_j (.sel(n_9), .in1(A[13]), .in2(), .i1(), .i2(), 
      .out1(sum[13]), .Carry(n_10));
   mux__15_197 muxx_14_muxx_j (.sel(n_10), .in1(A[14]), .in2(), .i1(), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__15_194 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__15_190(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_187(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_1 (.A(in1), .B(in2), .ZN(S));
endmodule

module FullAdder__15_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in2), .B(in1), .Z(S));
endmodule

module FullAdder__15_183(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_177(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_138(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_135(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_132(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_129(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_126(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_123(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_120(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_117(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_114(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_111(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_108(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_105(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__15_102(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__15_99(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_96(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_93(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_90(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_87(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_84(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_81(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__15_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_1_0 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module Addition1__15_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire S;
   wire Carry;

   FullAdder__15_190 FA0 (.in1(A[0]), .in2(B[0]), .Ci(), .S(sum[0]), .Co(n_0));
   FullAdder__15_187 FA_15_FA1_i (.in1(A[15]), .in2(B[15]), .Ci(), .S(S), .Co());
   FullAdder__15_185 FA_15_FA0_i (.in1(A[15]), .in2(B[15]), .Ci(), .S(n_2), 
      .Co());
   FullAdder__15_183 FA_14_FA1_i (.in1(A[14]), .in2(B[14]), .Ci(), .S(n_4), 
      .Co(n_3));
   FullAdder__15_180 FA_14_FA0_i (.in1(A[14]), .in2(B[14]), .Ci(), .S(n_6), 
      .Co(n_5));
   FullAdder__15_177 FA_13_FA1_i (.in1(A[13]), .in2(B[13]), .Ci(), .S(n_8), 
      .Co(n_7));
   FullAdder__15_174 FA_13_FA0_i (.in1(A[13]), .in2(B[13]), .Ci(), .S(n_10), 
      .Co(n_9));
   FullAdder__15_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__15_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__15_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__15_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__15_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__15_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__15_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__15_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__15_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__15_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_30), 
      .Co(n_29));
   FullAdder__15_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(n_32), 
      .Co(n_31));
   FullAdder__15_138 FA_7_FA0_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(n_34), 
      .Co(n_33));
   FullAdder__15_135 FA_6_FA1_i (.in1(A[6]), .in2(B[6]), .Ci(), .S(n_36), 
      .Co(n_35));
   FullAdder__15_132 FA_6_FA0_i (.in1(A[6]), .in2(B[6]), .Ci(), .S(n_38), 
      .Co(n_37));
   FullAdder__15_129 FA_5_FA1_i (.in1(A[5]), .in2(B[5]), .Ci(), .S(n_40), 
      .Co(n_39));
   FullAdder__15_126 FA_5_FA0_i (.in1(A[5]), .in2(B[5]), .Ci(), .S(n_42), 
      .Co(n_41));
   FullAdder__15_123 FA_4_FA1_i (.in1(A[4]), .in2(B[4]), .Ci(), .S(n_44), 
      .Co(n_43));
   FullAdder__15_120 FA_4_FA0_i (.in1(A[4]), .in2(B[4]), .Ci(), .S(n_46), 
      .Co(n_45));
   FullAdder__15_117 FA_3_FA1_i (.in1(A[3]), .in2(B[3]), .Ci(), .S(n_48), 
      .Co(n_47));
   FullAdder__15_114 FA_3_FA0_i (.in1(A[3]), .in2(B[3]), .Ci(), .S(n_50), 
      .Co(n_49));
   FullAdder__15_111 FA_2_FA1_i (.in1(A[2]), .in2(B[2]), .Ci(), .S(n_52), 
      .Co(n_51));
   FullAdder__15_108 FA_2_FA0_i (.in1(A[2]), .in2(B[2]), .Ci(), .S(n_54), 
      .Co(n_53));
   FullAdder__15_105 FA_1_FA1_i (.in1(A[1]), .in2(B[1]), .Ci(), .S(n_56), 
      .Co(n_55));
   FullAdder__15_102 FA_1_FA0_i (.in1(A[1]), .in2(B[1]), .Ci(), .S(n_58), 
      .Co(n_57));
   mux__15_99 muxx_1_muxx_j (.sel(n_0), .in1(n_58), .in2(n_56), .i1(n_57), 
      .i2(n_55), .out1(sum[1]), .Carry(n_59));
   mux__15_96 muxx_2_muxx_j (.sel(n_59), .in1(n_54), .in2(n_52), .i1(n_53), 
      .i2(n_51), .out1(sum[2]), .Carry(n_60));
   mux__15_93 muxx_3_muxx_j (.sel(n_60), .in1(n_50), .in2(n_48), .i1(n_49), 
      .i2(n_47), .out1(sum[3]), .Carry(n_61));
   mux__15_90 muxx_4_muxx_j (.sel(n_61), .in1(n_46), .in2(n_44), .i1(n_45), 
      .i2(n_43), .out1(sum[4]), .Carry(n_62));
   mux__15_87 muxx_5_muxx_j (.sel(n_62), .in1(n_42), .in2(n_40), .i1(n_41), 
      .i2(n_39), .out1(sum[5]), .Carry(n_63));
   mux__15_84 muxx_6_muxx_j (.sel(n_63), .in1(n_38), .in2(n_36), .i1(n_37), 
      .i2(n_35), .out1(sum[6]), .Carry(n_64));
   mux__15_81 muxx_7_muxx_j (.sel(n_64), .in1(n_34), .in2(n_32), .i1(n_33), 
      .i2(n_31), .out1(sum[7]), .Carry(n_65));
   mux__15_78 muxx_8_muxx_j (.sel(n_65), .in1(n_30), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_66));
   mux__15_75 muxx_9_muxx_j (.sel(n_66), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_67));
   mux__15_72 muxx_10_muxx_j (.sel(n_67), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_68));
   mux__15_69 muxx_11_muxx_j (.sel(n_68), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_69));
   mux__15_66 muxx_12_muxx_j (.sel(n_69), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_70));
   mux__15_63 muxx_13_muxx_j (.sel(n_70), .in1(n_10), .in2(n_8), .i1(n_9), 
      .i2(n_7), .out1(sum[13]), .Carry(n_1));
   mux__15_60 muxx_14_muxx_j (.sel(n_1), .in1(n_6), .in2(n_4), .i1(n_5), 
      .i2(n_3), .out1(sum[14]), .Carry(Carry));
   mux__15_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(S), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__15_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__15_191 u1 (.A(notplus), .B(firstVal), .Cin(), .sum({n_0, sum[14], 
      sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], sum[7], sum[6], sum[5], 
      sum[4], sum[3], sum[2], sum[1], sum[0]}), .overFlow());
   NOR4_X1 i_0_0 (.A1(sum[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(sum[6]), .A4(sum[5]), .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(sum[4]), .A2(sum[3]), .A3(sum[2]), .A4(sum[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_0 (.A(secondVal[0]), .ZN(notplus[0]));
   INV_X1 i_1_1 (.A(secondVal[1]), .ZN(notplus[1]));
   INV_X1 i_1_2 (.A(secondVal[2]), .ZN(notplus[2]));
   INV_X1 i_1_3 (.A(secondVal[3]), .ZN(notplus[3]));
   INV_X1 i_1_4 (.A(secondVal[4]), .ZN(notplus[4]));
   INV_X1 i_1_5 (.A(secondVal[5]), .ZN(notplus[5]));
   INV_X1 i_1_6 (.A(secondVal[6]), .ZN(notplus[6]));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
   INV_X1 i_1_13 (.A(secondVal[13]), .ZN(notplus[13]));
   INV_X1 i_1_14 (.A(secondVal[14]), .ZN(notplus[14]));
   INV_X1 i_1_15 (.A(secondVal[15]), .ZN(notplus[15]));
endmodule

module smallMux__15_53(loadAddress, CurrentCount, start, universalReset, 
      innerDone, continue, load, address);
   input [15:0]loadAddress;
   input [15:0]CurrentCount;
   input [15:0]start;
   input universalReset;
   input innerDone;
   input continue;
   input load;
   output [15:0]address;

   wire n_0_0;
   wire n_0_1;

   AND2_X1 i_0_0 (.A1(CurrentCount[0]), .A2(n_0_0), .ZN(address[0]));
   AND2_X1 i_0_1 (.A1(CurrentCount[1]), .A2(n_0_0), .ZN(address[1]));
   AND2_X1 i_0_2 (.A1(CurrentCount[2]), .A2(n_0_0), .ZN(address[2]));
   AND2_X1 i_0_3 (.A1(CurrentCount[3]), .A2(n_0_0), .ZN(address[3]));
   AND2_X1 i_0_4 (.A1(CurrentCount[4]), .A2(n_0_0), .ZN(address[4]));
   AND2_X1 i_0_5 (.A1(CurrentCount[5]), .A2(n_0_0), .ZN(address[5]));
   AND2_X1 i_0_6 (.A1(CurrentCount[6]), .A2(n_0_0), .ZN(address[6]));
   AND2_X1 i_0_7 (.A1(CurrentCount[7]), .A2(n_0_0), .ZN(address[7]));
   AND2_X1 i_0_8 (.A1(CurrentCount[8]), .A2(n_0_0), .ZN(address[8]));
   AND2_X1 i_0_9 (.A1(CurrentCount[9]), .A2(n_0_0), .ZN(address[9]));
   AND2_X1 i_0_10 (.A1(CurrentCount[10]), .A2(n_0_0), .ZN(address[10]));
   AND2_X1 i_0_11 (.A1(CurrentCount[11]), .A2(n_0_0), .ZN(address[11]));
   AND2_X1 i_0_12 (.A1(CurrentCount[12]), .A2(n_0_0), .ZN(address[12]));
   AND2_X1 i_0_13 (.A1(CurrentCount[13]), .A2(n_0_0), .ZN(address[13]));
   AND2_X1 i_0_14 (.A1(CurrentCount[14]), .A2(n_0_0), .ZN(address[14]));
   AND2_X1 i_0_15 (.A1(CurrentCount[15]), .A2(n_0_0), .ZN(address[15]));
   NOR2_X1 i_0_16 (.A1(n_0_1), .A2(universalReset), .ZN(n_0_0));
   NAND2_X1 i_0_17 (.A1(continue), .A2(innerDone), .ZN(n_0_1));
endmodule

module reg__15_49(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counterMux__15_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(n_0_0), .A2(counter[0]), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(counter[1]), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(counter[2]), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(counter[3]), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(counter[4]), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(counter[5]), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(counter[6]), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(counter[7]), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(counter[8]), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(counter[9]), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(counter[10]), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(counter[11]), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(counter[12]), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(counter[13]), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(counter[14]), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(counter[15]), .ZN(result[15]));
   INV_X1 i_0_16 (.A(universalReset), .ZN(n_0_0));
endmodule

module reg__15_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module flipflop__15_6(D, load, Clk, Q, rst);
   input D;
   input load;
   input Clk;
   output Q;
   input rst;

   DFFR_X1 Q_reg (.D(D), .RN(n_1), .CK(n_0), .Q(Q), .QN());
   INV_X1 i_0_0 (.A(Clk), .ZN(n_0));
   INV_X1 i_1_0 (.A(rst), .ZN(n_1));
endmodule

module counter__14_425(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]plus;
   wire [15:0]newStart;
   wire [15:0]init;
   wire [15:0]muxOut;
   wire n_0_1;
   wire n_0_0;
   wire activate;
   wire n_0_2;
   wire ffIN;
   wire setNewstart;

   Addition1__15_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   Addition1__15_328 u0 (.A({init[15], init[14], init[13], init[12], init[11], 
      init[10], init[9], init[8], init[7], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, 
      uc_6}), .B({uc_7, uc_8, uc_9, offset[12], offset[11], offset[10], 
      offset[9], offset[8], offset[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16}), .Cin(), .sum({plus[15], plus[14], plus[13], plus[12], plus[11], 
      plus[10], plus[9], plus[8], plus[7], uc_17, uc_18, uc_19, uc_20, uc_21, 
      uc_22, uc_23}), .overFlow());
   comparator__15_192 compare (.firstVal(dataOut), .secondVal({plus[15], 
      plus[14], plus[13], plus[12], plus[11], plus[10], plus[9], plus[8], 
      plus[7], init[6], init[5], init[4], init[3], init[2], init[1], init[0]}), 
      .done(done), .firstBigger(), .firstSmaller());
   smallMux__15_53 smallMux (.loadAddress(), .CurrentCount(dataOut), .start(), 
      .universalReset(universalReset), .innerDone(done), .continue(continue), 
      .load(), .address(newStart));
   reg__15_49 initialAdress (.D(newStart), .load(setNewstart), .Clk(CLK), 
      .Q(init), .rst(universalReset));
   counterMux__15_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(), .universalReset(universalReset), .continue(), 
      .result(muxOut));
   reg__15_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   flipflop__15_6 ff (.D(ffIN), .load(), .Clk(CLK), .Q(NFN), .rst(universalReset));
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(done), .ZN(n_0_1));
   INV_X1 i_0_1 (.A(enable), .ZN(n_0_0));
   OR2_X1 i_0_2 (.A1(n_0_1), .A2(universalReset), .ZN(activate));
   AND2_X1 i_0_3 (.A1(done), .A2(continue), .ZN(n_0_2));
   OR2_X1 i_0_4 (.A1(NFN), .A2(n_0_2), .ZN(ffIN));
   OR2_X1 i_0_5 (.A1(n_0_2), .A2(universalReset), .ZN(setNewstart));
endmodule

module FullAdder__17_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__17_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__17_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__17_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__17_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__17_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__17_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__17_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__17_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__17_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__17_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__17_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__17_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__17_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__17_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__17_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__17_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__17_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__17_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__17_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__17_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__17_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__17_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__17_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__17_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__17_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__17_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__17_185 FA_15_FA0_i (.in1(), .in2(B[15]), .Ci(), .S(n_2), .Co());
   FullAdder__17_180 FA_14_FA0_i (.in1(), .in2(B[14]), .Ci(), .S(n_6), .Co());
   FullAdder__17_174 FA_13_FA0_i (.in1(), .in2(B[13]), .Ci(), .S(n_10), .Co());
   FullAdder__17_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__17_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__17_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__17_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__17_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__17_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__17_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__17_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__17_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__17_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_0), 
      .Co(n_29));
   FullAdder__17_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_1));
   mux__17_78 muxx_8_muxx_j (.sel(n_1), .in1(n_0), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_3));
   mux__17_75 muxx_9_muxx_j (.sel(n_3), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_4));
   mux__17_72 muxx_10_muxx_j (.sel(n_4), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_5));
   mux__17_69 muxx_11_muxx_j (.sel(n_5), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_7));
   mux__17_66 muxx_12_muxx_j (.sel(n_7), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_8));
   mux__17_63 muxx_13_muxx_j (.sel(n_8), .in1(n_10), .in2(), .i1(B[13]), .i2(), 
      .out1(sum[13]), .Carry(n_9));
   mux__17_60 muxx_14_muxx_j (.sel(n_9), .in1(n_6), .in2(), .i1(B[14]), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__17_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__17_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__17_191 u1 (.A({uc_0, uc_1, uc_2, notplus[12], notplus[11], 
      notplus[10], notplus[9], notplus[8], notplus[7], uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9}), .B({firstVal[15], firstVal[14], firstVal[13], 
      firstVal[12], firstVal[11], firstVal[10], firstVal[9], firstVal[8], 
      firstVal[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16}), .Cin(), 
      .sum({n_0, sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
      sum[7], uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23}), .overFlow());
   NOR4_X1 i_0_0 (.A1(firstVal[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), 
      .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(firstVal[6]), .A4(firstVal[5]), 
      .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(firstVal[4]), .A2(firstVal[3]), .A3(firstVal[2]), .A4(
      firstVal[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
endmodule

module counterMux__17_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(counter[0]), .A2(n_0_0), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(counter[1]), .A2(n_0_0), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(counter[2]), .A2(n_0_0), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(counter[3]), .A2(n_0_0), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(counter[4]), .A2(n_0_0), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(counter[5]), .A2(n_0_0), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(counter[6]), .A2(n_0_0), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(counter[7]), .A2(n_0_0), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(counter[8]), .A2(n_0_0), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(counter[9]), .A2(n_0_0), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(counter[10]), .A2(n_0_0), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(counter[11]), .A2(n_0_0), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(counter[12]), .A2(n_0_0), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(counter[13]), .A2(n_0_0), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(counter[14]), .A2(n_0_0), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(counter[15]), .A2(n_0_0), .ZN(result[15]));
   NOR2_X1 i_0_16 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
endmodule

module reg__17_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__16_425(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]muxOut;
   wire activate;
   wire n_0_0;
   wire n_0_1;

   Addition1__17_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   comparator__17_192 compare (.firstVal(dataOut), .secondVal({uc_0, uc_1, uc_2, 
      offset[12], offset[11], offset[10], offset[9], offset[8], offset[7], uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .done(n_0), .firstBigger(), 
      .firstSmaller());
   counterMux__17_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(reset), .universalReset(universalReset), 
      .continue(), .result(muxOut));
   reg__17_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0), .ZN(activate));
   NOR2_X1 i_0_1 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(enable), .ZN(n_0_1));
endmodule

module FullAdder__17_423__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__17_392__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_389__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_386__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_383__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_380__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_377__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_374__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_371__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_368__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_365__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_362__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_359__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_356__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_353__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__17_350__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__17_424__1(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__17_423__1 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__17_392__1 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__17_389__1 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__17_386__1 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__17_383__1 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__17_380__1 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__17_377__1 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__17_374__1 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__17_371__1 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__17_368__1 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__17_365__1 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__17_362__1 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__17_359__1 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__17_356__1 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__17_353__1 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__17_350__1 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__17_185__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__17_180__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__17_174__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__17_171__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_168__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_165__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_162__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_159__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_156__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_153__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_150__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_147__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_144__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__17_141__1(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__17_78__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_75__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_72__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_69__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_66__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__17_63__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__17_60__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__17_57__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__17_191__1(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__17_185__1 FA_15_FA0_i (.in1(), .in2(B[15]), .Ci(), .S(n_2), .Co());
   FullAdder__17_180__1 FA_14_FA0_i (.in1(), .in2(B[14]), .Ci(), .S(n_6), .Co());
   FullAdder__17_174__1 FA_13_FA0_i (.in1(), .in2(B[13]), .Ci(), .S(n_10), .Co());
   FullAdder__17_171__1 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__17_168__1 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__17_165__1 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__17_162__1 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__17_159__1 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__17_156__1 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__17_153__1 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__17_150__1 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__17_147__1 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__17_144__1 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_0), 
      .Co(n_29));
   FullAdder__17_141__1 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_1));
   mux__17_78__1 muxx_8_muxx_j (.sel(n_1), .in1(n_0), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_3));
   mux__17_75__1 muxx_9_muxx_j (.sel(n_3), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_4));
   mux__17_72__1 muxx_10_muxx_j (.sel(n_4), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_5));
   mux__17_69__1 muxx_11_muxx_j (.sel(n_5), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_7));
   mux__17_66__1 muxx_12_muxx_j (.sel(n_7), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_8));
   mux__17_63__1 muxx_13_muxx_j (.sel(n_8), .in1(n_10), .in2(), .i1(B[13]), 
      .i2(), .out1(sum[13]), .Carry(n_9));
   mux__17_60__1 muxx_14_muxx_j (.sel(n_9), .in1(n_6), .in2(), .i1(B[14]), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__17_57__1 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__17_192__1(firstVal, secondVal, done, firstBigger, 
      firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__17_191__1 u1 (.A({uc_0, uc_1, uc_2, notplus[12], notplus[11], 
      notplus[10], notplus[9], notplus[8], notplus[7], uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9}), .B({firstVal[15], firstVal[14], firstVal[13], 
      firstVal[12], firstVal[11], firstVal[10], firstVal[9], firstVal[8], 
      firstVal[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16}), .Cin(), 
      .sum({n_0, sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
      sum[7], uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23}), .overFlow());
   NOR4_X1 i_0_0 (.A1(firstVal[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), 
      .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(firstVal[6]), .A4(firstVal[5]), 
      .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(firstVal[4]), .A2(firstVal[3]), .A3(firstVal[2]), .A4(
      firstVal[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
endmodule

module counterMux__17_29__1(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(counter[0]), .A2(n_0_0), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(counter[1]), .A2(n_0_0), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(counter[2]), .A2(n_0_0), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(counter[3]), .A2(n_0_0), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(counter[4]), .A2(n_0_0), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(counter[5]), .A2(n_0_0), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(counter[6]), .A2(n_0_0), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(counter[7]), .A2(n_0_0), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(counter[8]), .A2(n_0_0), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(counter[9]), .A2(n_0_0), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(counter[10]), .A2(n_0_0), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(counter[11]), .A2(n_0_0), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(counter[12]), .A2(n_0_0), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(counter[13]), .A2(n_0_0), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(counter[14]), .A2(n_0_0), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(counter[15]), .A2(n_0_0), .ZN(result[15]));
   NOR2_X1 i_0_16 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
endmodule

module reg__17_26__1(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__16_425__1(dataIn, offset, load, enable, CLK, reset, 
      universalReset, continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]muxOut;
   wire activate;
   wire n_0_0;
   wire n_0_1;

   Addition1__17_424__1 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   comparator__17_192__1 compare (.firstVal(dataOut), .secondVal({uc_0, uc_1, 
      uc_2, offset[12], offset[11], offset[10], offset[9], offset[8], offset[7], 
      uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .done(n_0), .firstBigger(), 
      .firstSmaller());
   counterMux__17_29__1 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(reset), .universalReset(universalReset), 
      .continue(), .result(muxOut));
   reg__17_26__1 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0), .ZN(activate));
   NOR2_X1 i_0_1 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(enable), .ZN(n_0_1));
endmodule

module FullAdder__18_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__18_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__18_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__18_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__18_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__18_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__18_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__18_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__18_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__18_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__18_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__18_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__18_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__18_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__18_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__18_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__18_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__18_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__18_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__18_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__18_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__18_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__18_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__18_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__18_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__18_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__18_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__18_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__18_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__18_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__18_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__18_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__18_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__18_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__18_185 FA_15_FA0_i (.in1(), .in2(B[15]), .Ci(), .S(n_2), .Co());
   FullAdder__18_180 FA_14_FA0_i (.in1(), .in2(B[14]), .Ci(), .S(n_6), .Co());
   FullAdder__18_174 FA_13_FA0_i (.in1(), .in2(B[13]), .Ci(), .S(n_10), .Co());
   FullAdder__18_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__18_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__18_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__18_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__18_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__18_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__18_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__18_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__18_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__18_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_0), 
      .Co(n_29));
   FullAdder__18_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_1));
   mux__18_78 muxx_8_muxx_j (.sel(n_1), .in1(n_0), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_3));
   mux__18_75 muxx_9_muxx_j (.sel(n_3), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_4));
   mux__18_72 muxx_10_muxx_j (.sel(n_4), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_5));
   mux__18_69 muxx_11_muxx_j (.sel(n_5), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_7));
   mux__18_66 muxx_12_muxx_j (.sel(n_7), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_8));
   mux__18_63 muxx_13_muxx_j (.sel(n_8), .in1(n_10), .in2(), .i1(B[13]), .i2(), 
      .out1(sum[13]), .Carry(n_9));
   mux__18_60 muxx_14_muxx_j (.sel(n_9), .in1(n_6), .in2(), .i1(B[14]), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__18_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__18_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__18_191 u1 (.A({uc_0, uc_1, uc_2, notplus[12], notplus[11], 
      notplus[10], notplus[9], notplus[8], notplus[7], uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9}), .B({firstVal[15], firstVal[14], firstVal[13], 
      firstVal[12], firstVal[11], firstVal[10], firstVal[9], firstVal[8], 
      firstVal[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16}), .Cin(), 
      .sum({n_0, sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
      sum[7], uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23}), .overFlow());
   NOR4_X1 i_0_0 (.A1(firstVal[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), 
      .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(firstVal[6]), .A4(firstVal[5]), 
      .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(firstVal[4]), .A2(firstVal[3]), .A3(firstVal[2]), .A4(
      firstVal[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
endmodule

module counterMux__18_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(counter[0]), .A2(n_0_0), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(counter[1]), .A2(n_0_0), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(counter[2]), .A2(n_0_0), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(counter[3]), .A2(n_0_0), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(counter[4]), .A2(n_0_0), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(counter[5]), .A2(n_0_0), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(counter[6]), .A2(n_0_0), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(counter[7]), .A2(n_0_0), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(counter[8]), .A2(n_0_0), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(counter[9]), .A2(n_0_0), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(counter[10]), .A2(n_0_0), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(counter[11]), .A2(n_0_0), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(counter[12]), .A2(n_0_0), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(counter[13]), .A2(n_0_0), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(counter[14]), .A2(n_0_0), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(counter[15]), .A2(n_0_0), .ZN(result[15]));
   NOR2_X1 i_0_16 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
endmodule

module reg__18_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__17_425(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]muxOut;
   wire activate;
   wire n_0_0;
   wire n_0_1;

   Addition1__18_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   comparator__18_192 compare (.firstVal(dataOut), .secondVal({uc_0, uc_1, uc_2, 
      offset[12], offset[11], offset[10], offset[9], offset[8], offset[7], uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .done(n_0), .firstBigger(), 
      .firstSmaller());
   counterMux__18_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(reset), .universalReset(universalReset), 
      .continue(), .result(muxOut));
   reg__18_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0), .ZN(activate));
   NOR2_X1 i_0_1 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(enable), .ZN(n_0_1));
endmodule

module FullAdder__19_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__19_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__19_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__19_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__19_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__19_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__19_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__19_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__19_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__19_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__19_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__19_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__19_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__19_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__19_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__19_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__19_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__19_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__19_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__19_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__19_308(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_305(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_302(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_299(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_296(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_293(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_290(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_287(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_284(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_281(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_275(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__19_215(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_212(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_209(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_206(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_203(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_200(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_0_0 (.A(in1), .B(sel), .Z(out1));
   AND2_X1 i_0_1 (.A1(sel), .A2(in1), .ZN(Carry));
endmodule

module mux__19_197(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_0_0 (.A(in1), .B(sel), .Z(out1));
   AND2_X1 i_0_1 (.A1(sel), .A2(in1), .ZN(Carry));
endmodule

module mux__19_194(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__19_328(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__19_308 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__19_305 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__19_302 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__19_299 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__19_296 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__19_293 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__19_290 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__19_287 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__19_284 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_1), 
      .Co(n_0));
   FullAdder__19_281 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_3), 
      .Co(n_2));
   FullAdder__19_275 FA_7_FA0_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_4));
   mux__19_215 muxx_8_muxx_j (.sel(n_4), .in1(n_3), .in2(n_1), .i1(n_2), 
      .i2(n_0), .out1(sum[8]), .Carry(n_5));
   mux__19_212 muxx_9_muxx_j (.sel(n_5), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_6));
   mux__19_209 muxx_10_muxx_j (.sel(n_6), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_7));
   mux__19_206 muxx_11_muxx_j (.sel(n_7), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_8));
   mux__19_203 muxx_12_muxx_j (.sel(n_8), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_9));
   mux__19_200 muxx_13_muxx_j (.sel(n_9), .in1(A[13]), .in2(), .i1(), .i2(), 
      .out1(sum[13]), .Carry(n_10));
   mux__19_197 muxx_14_muxx_j (.sel(n_10), .in1(A[14]), .in2(), .i1(), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__19_194 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__19_190(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_187(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_1 (.A(in1), .B(in2), .ZN(S));
endmodule

module FullAdder__19_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in2), .B(in1), .Z(S));
endmodule

module FullAdder__19_183(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_177(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_138(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_135(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_132(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_129(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_126(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_123(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_120(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_117(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_114(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_111(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_108(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_105(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__19_102(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__19_99(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_96(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_93(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_90(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_87(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_84(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_81(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__19_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_1_0 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module Addition1__19_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire S;
   wire Carry;

   FullAdder__19_190 FA0 (.in1(A[0]), .in2(B[0]), .Ci(), .S(sum[0]), .Co(n_0));
   FullAdder__19_187 FA_15_FA1_i (.in1(A[15]), .in2(B[15]), .Ci(), .S(S), .Co());
   FullAdder__19_185 FA_15_FA0_i (.in1(A[15]), .in2(B[15]), .Ci(), .S(n_2), 
      .Co());
   FullAdder__19_183 FA_14_FA1_i (.in1(A[14]), .in2(B[14]), .Ci(), .S(n_4), 
      .Co(n_3));
   FullAdder__19_180 FA_14_FA0_i (.in1(A[14]), .in2(B[14]), .Ci(), .S(n_6), 
      .Co(n_5));
   FullAdder__19_177 FA_13_FA1_i (.in1(A[13]), .in2(B[13]), .Ci(), .S(n_8), 
      .Co(n_7));
   FullAdder__19_174 FA_13_FA0_i (.in1(A[13]), .in2(B[13]), .Ci(), .S(n_10), 
      .Co(n_9));
   FullAdder__19_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__19_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__19_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__19_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__19_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__19_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__19_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__19_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__19_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__19_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_30), 
      .Co(n_29));
   FullAdder__19_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(n_32), 
      .Co(n_31));
   FullAdder__19_138 FA_7_FA0_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(n_34), 
      .Co(n_33));
   FullAdder__19_135 FA_6_FA1_i (.in1(A[6]), .in2(B[6]), .Ci(), .S(n_36), 
      .Co(n_35));
   FullAdder__19_132 FA_6_FA0_i (.in1(A[6]), .in2(B[6]), .Ci(), .S(n_38), 
      .Co(n_37));
   FullAdder__19_129 FA_5_FA1_i (.in1(A[5]), .in2(B[5]), .Ci(), .S(n_40), 
      .Co(n_39));
   FullAdder__19_126 FA_5_FA0_i (.in1(A[5]), .in2(B[5]), .Ci(), .S(n_42), 
      .Co(n_41));
   FullAdder__19_123 FA_4_FA1_i (.in1(A[4]), .in2(B[4]), .Ci(), .S(n_44), 
      .Co(n_43));
   FullAdder__19_120 FA_4_FA0_i (.in1(A[4]), .in2(B[4]), .Ci(), .S(n_46), 
      .Co(n_45));
   FullAdder__19_117 FA_3_FA1_i (.in1(A[3]), .in2(B[3]), .Ci(), .S(n_48), 
      .Co(n_47));
   FullAdder__19_114 FA_3_FA0_i (.in1(A[3]), .in2(B[3]), .Ci(), .S(n_50), 
      .Co(n_49));
   FullAdder__19_111 FA_2_FA1_i (.in1(A[2]), .in2(B[2]), .Ci(), .S(n_52), 
      .Co(n_51));
   FullAdder__19_108 FA_2_FA0_i (.in1(A[2]), .in2(B[2]), .Ci(), .S(n_54), 
      .Co(n_53));
   FullAdder__19_105 FA_1_FA1_i (.in1(A[1]), .in2(B[1]), .Ci(), .S(n_56), 
      .Co(n_55));
   FullAdder__19_102 FA_1_FA0_i (.in1(A[1]), .in2(B[1]), .Ci(), .S(n_58), 
      .Co(n_57));
   mux__19_99 muxx_1_muxx_j (.sel(n_0), .in1(n_58), .in2(n_56), .i1(n_57), 
      .i2(n_55), .out1(sum[1]), .Carry(n_59));
   mux__19_96 muxx_2_muxx_j (.sel(n_59), .in1(n_54), .in2(n_52), .i1(n_53), 
      .i2(n_51), .out1(sum[2]), .Carry(n_60));
   mux__19_93 muxx_3_muxx_j (.sel(n_60), .in1(n_50), .in2(n_48), .i1(n_49), 
      .i2(n_47), .out1(sum[3]), .Carry(n_61));
   mux__19_90 muxx_4_muxx_j (.sel(n_61), .in1(n_46), .in2(n_44), .i1(n_45), 
      .i2(n_43), .out1(sum[4]), .Carry(n_62));
   mux__19_87 muxx_5_muxx_j (.sel(n_62), .in1(n_42), .in2(n_40), .i1(n_41), 
      .i2(n_39), .out1(sum[5]), .Carry(n_63));
   mux__19_84 muxx_6_muxx_j (.sel(n_63), .in1(n_38), .in2(n_36), .i1(n_37), 
      .i2(n_35), .out1(sum[6]), .Carry(n_64));
   mux__19_81 muxx_7_muxx_j (.sel(n_64), .in1(n_34), .in2(n_32), .i1(n_33), 
      .i2(n_31), .out1(sum[7]), .Carry(n_65));
   mux__19_78 muxx_8_muxx_j (.sel(n_65), .in1(n_30), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_66));
   mux__19_75 muxx_9_muxx_j (.sel(n_66), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_67));
   mux__19_72 muxx_10_muxx_j (.sel(n_67), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_68));
   mux__19_69 muxx_11_muxx_j (.sel(n_68), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_69));
   mux__19_66 muxx_12_muxx_j (.sel(n_69), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_70));
   mux__19_63 muxx_13_muxx_j (.sel(n_70), .in1(n_10), .in2(n_8), .i1(n_9), 
      .i2(n_7), .out1(sum[13]), .Carry(n_1));
   mux__19_60 muxx_14_muxx_j (.sel(n_1), .in1(n_6), .in2(n_4), .i1(n_5), 
      .i2(n_3), .out1(sum[14]), .Carry(Carry));
   mux__19_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(S), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__19_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__19_191 u1 (.A(notplus), .B(firstVal), .Cin(), .sum({n_0, sum[14], 
      sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], sum[7], sum[6], sum[5], 
      sum[4], sum[3], sum[2], sum[1], sum[0]}), .overFlow());
   NOR4_X1 i_0_0 (.A1(sum[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(sum[6]), .A4(sum[5]), .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(sum[4]), .A2(sum[3]), .A3(sum[2]), .A4(sum[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_0 (.A(secondVal[0]), .ZN(notplus[0]));
   INV_X1 i_1_1 (.A(secondVal[1]), .ZN(notplus[1]));
   INV_X1 i_1_2 (.A(secondVal[2]), .ZN(notplus[2]));
   INV_X1 i_1_3 (.A(secondVal[3]), .ZN(notplus[3]));
   INV_X1 i_1_4 (.A(secondVal[4]), .ZN(notplus[4]));
   INV_X1 i_1_5 (.A(secondVal[5]), .ZN(notplus[5]));
   INV_X1 i_1_6 (.A(secondVal[6]), .ZN(notplus[6]));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
   INV_X1 i_1_13 (.A(secondVal[13]), .ZN(notplus[13]));
   INV_X1 i_1_14 (.A(secondVal[14]), .ZN(notplus[14]));
   INV_X1 i_1_15 (.A(secondVal[15]), .ZN(notplus[15]));
endmodule

module smallMux__19_53(loadAddress, CurrentCount, start, universalReset, 
      innerDone, continue, load, address);
   input [15:0]loadAddress;
   input [15:0]CurrentCount;
   input [15:0]start;
   input universalReset;
   input innerDone;
   input continue;
   input load;
   output [15:0]address;

   wire n_0_0;
   wire n_0_1;

   AND2_X1 i_0_0 (.A1(CurrentCount[0]), .A2(n_0_0), .ZN(address[0]));
   AND2_X1 i_0_1 (.A1(CurrentCount[1]), .A2(n_0_0), .ZN(address[1]));
   AND2_X1 i_0_2 (.A1(CurrentCount[2]), .A2(n_0_0), .ZN(address[2]));
   AND2_X1 i_0_3 (.A1(CurrentCount[3]), .A2(n_0_0), .ZN(address[3]));
   AND2_X1 i_0_4 (.A1(CurrentCount[4]), .A2(n_0_0), .ZN(address[4]));
   AND2_X1 i_0_5 (.A1(CurrentCount[5]), .A2(n_0_0), .ZN(address[5]));
   AND2_X1 i_0_6 (.A1(CurrentCount[6]), .A2(n_0_0), .ZN(address[6]));
   AND2_X1 i_0_7 (.A1(CurrentCount[7]), .A2(n_0_0), .ZN(address[7]));
   AND2_X1 i_0_8 (.A1(CurrentCount[8]), .A2(n_0_0), .ZN(address[8]));
   AND2_X1 i_0_9 (.A1(CurrentCount[9]), .A2(n_0_0), .ZN(address[9]));
   AND2_X1 i_0_10 (.A1(CurrentCount[10]), .A2(n_0_0), .ZN(address[10]));
   AND2_X1 i_0_11 (.A1(CurrentCount[11]), .A2(n_0_0), .ZN(address[11]));
   AND2_X1 i_0_12 (.A1(CurrentCount[12]), .A2(n_0_0), .ZN(address[12]));
   AND2_X1 i_0_13 (.A1(CurrentCount[13]), .A2(n_0_0), .ZN(address[13]));
   AND2_X1 i_0_14 (.A1(CurrentCount[14]), .A2(n_0_0), .ZN(address[14]));
   AND2_X1 i_0_15 (.A1(CurrentCount[15]), .A2(n_0_0), .ZN(address[15]));
   NOR2_X1 i_0_16 (.A1(n_0_1), .A2(universalReset), .ZN(n_0_0));
   NAND2_X1 i_0_17 (.A1(continue), .A2(innerDone), .ZN(n_0_1));
endmodule

module reg__19_49(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counterMux__19_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(n_0_0), .A2(counter[0]), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(counter[1]), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(counter[2]), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(counter[3]), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(counter[4]), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(counter[5]), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(counter[6]), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(counter[7]), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(counter[8]), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(counter[9]), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(counter[10]), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(counter[11]), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(counter[12]), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(counter[13]), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(counter[14]), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(counter[15]), .ZN(result[15]));
   INV_X1 i_0_16 (.A(universalReset), .ZN(n_0_0));
endmodule

module reg__19_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__18_425(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]plus;
   wire [15:0]newStart;
   wire [15:0]init;
   wire [15:0]muxOut;
   wire setNewstart;
   wire n_0_0;
   wire activate;
   wire n_0_1;
   wire n_0_2;

   Addition1__19_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   Addition1__19_328 u0 (.A({init[15], init[14], init[13], init[12], init[11], 
      init[10], init[9], init[8], init[7], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, 
      uc_6}), .B({uc_7, uc_8, uc_9, offset[12], offset[11], offset[10], 
      offset[9], offset[8], offset[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16}), .Cin(), .sum({plus[15], plus[14], plus[13], plus[12], plus[11], 
      plus[10], plus[9], plus[8], plus[7], uc_17, uc_18, uc_19, uc_20, uc_21, 
      uc_22, uc_23}), .overFlow());
   comparator__19_192 compare (.firstVal(dataOut), .secondVal({plus[15], 
      plus[14], plus[13], plus[12], plus[11], plus[10], plus[9], plus[8], 
      plus[7], init[6], init[5], init[4], init[3], init[2], init[1], init[0]}), 
      .done(n_0), .firstBigger(), .firstSmaller());
   smallMux__19_53 smallMux (.loadAddress(), .CurrentCount(dataOut), .start(), 
      .universalReset(universalReset), .innerDone(n_0), .continue(continue), 
      .load(), .address(newStart));
   reg__19_49 initialAdress (.D(newStart), .load(setNewstart), .Clk(CLK), 
      .Q(init), .rst(universalReset));
   counterMux__19_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(), .universalReset(universalReset), .continue(), 
      .result(muxOut));
   reg__19_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   INV_X1 i_0_0 (.A(n_0_0), .ZN(setNewstart));
   AOI21_X1 i_0_1 (.A(universalReset), .B1(n_0), .B2(continue), .ZN(n_0_0));
   OAI21_X1 i_0_2 (.A(n_0_2), .B1(n_0_1), .B2(n_0), .ZN(activate));
   INV_X1 i_0_3 (.A(enable), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(universalReset), .ZN(n_0_2));
endmodule

module FullAdder__20_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__20_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__20_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__20_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__20_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__20_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__20_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__20_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__20_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__20_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__20_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__20_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__20_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__20_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__20_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__20_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__20_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__20_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__20_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__20_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__20_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__20_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__20_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__20_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__20_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__20_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__20_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__20_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__20_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__20_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__20_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__20_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__20_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__20_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__20_185 FA_15_FA0_i (.in1(), .in2(B[15]), .Ci(), .S(n_2), .Co());
   FullAdder__20_180 FA_14_FA0_i (.in1(), .in2(B[14]), .Ci(), .S(n_6), .Co());
   FullAdder__20_174 FA_13_FA0_i (.in1(), .in2(B[13]), .Ci(), .S(n_10), .Co());
   FullAdder__20_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__20_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__20_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__20_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__20_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__20_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__20_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__20_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__20_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__20_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_0), 
      .Co(n_29));
   FullAdder__20_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_1));
   mux__20_78 muxx_8_muxx_j (.sel(n_1), .in1(n_0), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_3));
   mux__20_75 muxx_9_muxx_j (.sel(n_3), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_4));
   mux__20_72 muxx_10_muxx_j (.sel(n_4), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_5));
   mux__20_69 muxx_11_muxx_j (.sel(n_5), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_7));
   mux__20_66 muxx_12_muxx_j (.sel(n_7), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_8));
   mux__20_63 muxx_13_muxx_j (.sel(n_8), .in1(n_10), .in2(), .i1(B[13]), .i2(), 
      .out1(sum[13]), .Carry(n_9));
   mux__20_60 muxx_14_muxx_j (.sel(n_9), .in1(n_6), .in2(), .i1(B[14]), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__20_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__20_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__20_191 u1 (.A({uc_0, uc_1, uc_2, notplus[12], notplus[11], 
      notplus[10], notplus[9], notplus[8], notplus[7], uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9}), .B({firstVal[15], firstVal[14], firstVal[13], 
      firstVal[12], firstVal[11], firstVal[10], firstVal[9], firstVal[8], 
      firstVal[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16}), .Cin(), 
      .sum({n_0, sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
      sum[7], uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23}), .overFlow());
   NOR4_X1 i_0_0 (.A1(firstVal[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), 
      .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(firstVal[6]), .A4(firstVal[5]), 
      .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(firstVal[4]), .A2(firstVal[3]), .A3(firstVal[2]), .A4(
      firstVal[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
endmodule

module counterMux__20_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(counter[0]), .A2(n_0_0), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(counter[1]), .A2(n_0_0), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(counter[2]), .A2(n_0_0), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(counter[3]), .A2(n_0_0), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(counter[4]), .A2(n_0_0), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(counter[5]), .A2(n_0_0), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(counter[6]), .A2(n_0_0), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(counter[7]), .A2(n_0_0), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(counter[8]), .A2(n_0_0), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(counter[9]), .A2(n_0_0), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(counter[10]), .A2(n_0_0), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(counter[11]), .A2(n_0_0), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(counter[12]), .A2(n_0_0), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(counter[13]), .A2(n_0_0), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(counter[14]), .A2(n_0_0), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(counter[15]), .A2(n_0_0), .ZN(result[15]));
   NOR2_X1 i_0_16 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
endmodule

module reg__20_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__19_425(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]muxOut;
   wire activate;
   wire n_0_0;
   wire n_0_1;

   Addition1__20_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   comparator__20_192 compare (.firstVal(dataOut), .secondVal({uc_0, uc_1, uc_2, 
      offset[12], offset[11], offset[10], offset[9], offset[8], offset[7], uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .done(n_0), .firstBigger(), 
      .firstSmaller());
   counterMux__20_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(reset), .universalReset(universalReset), 
      .continue(), .result(muxOut));
   reg__20_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0), .ZN(activate));
   NOR2_X1 i_0_1 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(enable), .ZN(n_0_1));
endmodule

module FullAdder__21_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__21_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__21_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__21_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__21_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__21_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__21_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__21_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__21_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__21_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__21_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__21_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__21_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__21_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__21_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__21_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__21_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__21_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__21_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__21_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__21_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__21_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__21_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__21_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__21_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__21_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__21_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__21_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__21_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__21_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__21_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__21_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__21_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__21_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__21_185 FA_15_FA0_i (.in1(), .in2(B[15]), .Ci(), .S(n_2), .Co());
   FullAdder__21_180 FA_14_FA0_i (.in1(), .in2(B[14]), .Ci(), .S(n_6), .Co());
   FullAdder__21_174 FA_13_FA0_i (.in1(), .in2(B[13]), .Ci(), .S(n_10), .Co());
   FullAdder__21_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__21_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__21_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__21_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__21_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__21_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__21_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__21_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__21_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__21_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_0), 
      .Co(n_29));
   FullAdder__21_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_1));
   mux__21_78 muxx_8_muxx_j (.sel(n_1), .in1(n_0), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_3));
   mux__21_75 muxx_9_muxx_j (.sel(n_3), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_4));
   mux__21_72 muxx_10_muxx_j (.sel(n_4), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_5));
   mux__21_69 muxx_11_muxx_j (.sel(n_5), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_7));
   mux__21_66 muxx_12_muxx_j (.sel(n_7), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_8));
   mux__21_63 muxx_13_muxx_j (.sel(n_8), .in1(n_10), .in2(), .i1(B[13]), .i2(), 
      .out1(sum[13]), .Carry(n_9));
   mux__21_60 muxx_14_muxx_j (.sel(n_9), .in1(n_6), .in2(), .i1(B[14]), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__21_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__21_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__21_191 u1 (.A({uc_0, uc_1, uc_2, notplus[12], notplus[11], 
      notplus[10], notplus[9], notplus[8], notplus[7], uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9}), .B({firstVal[15], firstVal[14], firstVal[13], 
      firstVal[12], firstVal[11], firstVal[10], firstVal[9], firstVal[8], 
      firstVal[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16}), .Cin(), 
      .sum({n_0, sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
      sum[7], uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23}), .overFlow());
   NOR4_X1 i_0_0 (.A1(firstVal[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), 
      .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(firstVal[6]), .A4(firstVal[5]), 
      .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(firstVal[4]), .A2(firstVal[3]), .A3(firstVal[2]), .A4(
      firstVal[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
endmodule

module counterMux__21_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(counter[0]), .A2(n_0_0), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(counter[1]), .A2(n_0_0), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(counter[2]), .A2(n_0_0), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(counter[3]), .A2(n_0_0), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(counter[4]), .A2(n_0_0), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(counter[5]), .A2(n_0_0), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(counter[6]), .A2(n_0_0), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(counter[7]), .A2(n_0_0), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(counter[8]), .A2(n_0_0), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(counter[9]), .A2(n_0_0), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(counter[10]), .A2(n_0_0), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(counter[11]), .A2(n_0_0), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(counter[12]), .A2(n_0_0), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(counter[13]), .A2(n_0_0), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(counter[14]), .A2(n_0_0), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(counter[15]), .A2(n_0_0), .ZN(result[15]));
   NOR2_X1 i_0_16 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
endmodule

module reg__21_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__20_425(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]muxOut;
   wire activate;
   wire n_0_0;
   wire n_0_1;

   Addition1__21_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   comparator__21_192 compare (.firstVal(dataOut), .secondVal({uc_0, uc_1, uc_2, 
      offset[12], offset[11], offset[10], offset[9], offset[8], offset[7], uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .done(n_0), .firstBigger(), 
      .firstSmaller());
   counterMux__21_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(reset), .universalReset(universalReset), 
      .continue(), .result(muxOut));
   reg__21_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0), .ZN(activate));
   NOR2_X1 i_0_1 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(enable), .ZN(n_0_1));
endmodule

module FullAdder__22_423(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_2 (.A(in1), .ZN(S));
endmodule

module mux__22_392(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_389(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_386(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_383(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_380(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_377(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_374(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_371(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_368(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_365(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_362(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_359(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_356(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_353(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__22_350(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__22_424(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__22_423 FA0 (.in1(A[0]), .in2(), .Ci(), .S(sum[0]), .Co());
   mux__22_392 muxx_1_muxx_j (.sel(A[0]), .in1(), .in2(), .i1(), .i2(A[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__22_389 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(A[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__22_386 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(A[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__22_383 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(A[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__22_380 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(A[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__22_377 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(A[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__22_374 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(A[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__22_371 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(A[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__22_368 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(A[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__22_365 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(A[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__22_362 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(A[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__22_359 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(A[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__22_356 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(A[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__22_353 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(A[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__22_350 muxx_15_muxx_j (.sel(Carry), .in1(A[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module FullAdder__22_185(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__22_180(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__22_174(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   INV_X1 i_0_0 (.A(in2), .ZN(S));
endmodule

module FullAdder__22_171(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_168(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_165(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_162(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_159(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_156(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_153(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_150(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_147(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_144(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XOR2_X1 i_0_0 (.A(in1), .B(in2), .Z(S));
   AND2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module FullAdder__22_141(in1, in2, Ci, S, Co);
   input in1;
   input in2;
   input Ci;
   output S;
   output Co;

   XNOR2_X1 i_0_0 (.A(in2), .B(in1), .ZN(S));
   OR2_X1 i_0_1 (.A1(in2), .A2(in1), .ZN(Co));
endmodule

module mux__22_78(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__22_75(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__22_72(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__22_69(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__22_66(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   MUX2_X1 i_0_0 (.A(i1), .B(i2), .S(sel), .Z(Carry));
   MUX2_X1 i_0_1 (.A(in1), .B(in2), .S(sel), .Z(out1));
endmodule

module mux__22_63(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__22_60(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   OR2_X1 i_0_0 (.A1(sel), .A2(i1), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(in1), .B(sel), .Z(out1));
endmodule

module mux__22_57(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__22_191(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   FullAdder__22_185 FA_15_FA0_i (.in1(), .in2(B[15]), .Ci(), .S(n_2), .Co());
   FullAdder__22_180 FA_14_FA0_i (.in1(), .in2(B[14]), .Ci(), .S(n_6), .Co());
   FullAdder__22_174 FA_13_FA0_i (.in1(), .in2(B[13]), .Ci(), .S(n_10), .Co());
   FullAdder__22_171 FA_12_FA1_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_12), 
      .Co(n_11));
   FullAdder__22_168 FA_12_FA0_i (.in1(A[12]), .in2(B[12]), .Ci(), .S(n_14), 
      .Co(n_13));
   FullAdder__22_165 FA_11_FA1_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_16), 
      .Co(n_15));
   FullAdder__22_162 FA_11_FA0_i (.in1(A[11]), .in2(B[11]), .Ci(), .S(n_18), 
      .Co(n_17));
   FullAdder__22_159 FA_10_FA1_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_20), 
      .Co(n_19));
   FullAdder__22_156 FA_10_FA0_i (.in1(A[10]), .in2(B[10]), .Ci(), .S(n_22), 
      .Co(n_21));
   FullAdder__22_153 FA_9_FA1_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_24), 
      .Co(n_23));
   FullAdder__22_150 FA_9_FA0_i (.in1(A[9]), .in2(B[9]), .Ci(), .S(n_26), 
      .Co(n_25));
   FullAdder__22_147 FA_8_FA1_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_28), 
      .Co(n_27));
   FullAdder__22_144 FA_8_FA0_i (.in1(A[8]), .in2(B[8]), .Ci(), .S(n_0), 
      .Co(n_29));
   FullAdder__22_141 FA_7_FA1_i (.in1(A[7]), .in2(B[7]), .Ci(), .S(sum[7]), 
      .Co(n_1));
   mux__22_78 muxx_8_muxx_j (.sel(n_1), .in1(n_0), .in2(n_28), .i1(n_29), 
      .i2(n_27), .out1(sum[8]), .Carry(n_3));
   mux__22_75 muxx_9_muxx_j (.sel(n_3), .in1(n_26), .in2(n_24), .i1(n_25), 
      .i2(n_23), .out1(sum[9]), .Carry(n_4));
   mux__22_72 muxx_10_muxx_j (.sel(n_4), .in1(n_22), .in2(n_20), .i1(n_21), 
      .i2(n_19), .out1(sum[10]), .Carry(n_5));
   mux__22_69 muxx_11_muxx_j (.sel(n_5), .in1(n_18), .in2(n_16), .i1(n_17), 
      .i2(n_15), .out1(sum[11]), .Carry(n_7));
   mux__22_66 muxx_12_muxx_j (.sel(n_7), .in1(n_14), .in2(n_12), .i1(n_13), 
      .i2(n_11), .out1(sum[12]), .Carry(n_8));
   mux__22_63 muxx_13_muxx_j (.sel(n_8), .in1(n_10), .in2(), .i1(B[13]), .i2(), 
      .out1(sum[13]), .Carry(n_9));
   mux__22_60 muxx_14_muxx_j (.sel(n_9), .in1(n_6), .in2(), .i1(B[14]), .i2(), 
      .out1(sum[14]), .Carry(Carry));
   mux__22_57 muxx_15_muxx_j (.sel(Carry), .in1(n_2), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module comparator__22_192(firstVal, secondVal, done, firstBigger, firstSmaller);
   input [15:0]firstVal;
   input [15:0]secondVal;
   output done;
   output firstBigger;
   output firstSmaller;

   wire [15:0]sum;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire [15:0]notplus;

   Addition1__22_191 u1 (.A({uc_0, uc_1, uc_2, notplus[12], notplus[11], 
      notplus[10], notplus[9], notplus[8], notplus[7], uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9}), .B({firstVal[15], firstVal[14], firstVal[13], 
      firstVal[12], firstVal[11], firstVal[10], firstVal[9], firstVal[8], 
      firstVal[7], uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16}), .Cin(), 
      .sum({n_0, sum[14], sum[13], sum[12], sum[11], sum[10], sum[9], sum[8], 
      sum[7], uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23}), .overFlow());
   NOR4_X1 i_0_0 (.A1(firstVal[0]), .A2(n_0), .A3(sum[14]), .A4(sum[13]), 
      .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(sum[12]), .A2(sum[11]), .A3(sum[10]), .A4(sum[9]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(sum[8]), .A2(sum[7]), .A3(firstVal[6]), .A4(firstVal[5]), 
      .ZN(n_0_2));
   NOR4_X1 i_0_3 (.A1(firstVal[4]), .A2(firstVal[3]), .A3(firstVal[2]), .A4(
      firstVal[1]), .ZN(n_0_3));
   AND4_X1 i_0_4 (.A1(n_0_0), .A2(n_0_1), .A3(n_0_2), .A4(n_0_3), .ZN(done));
   INV_X1 i_1_7 (.A(secondVal[7]), .ZN(notplus[7]));
   INV_X1 i_1_8 (.A(secondVal[8]), .ZN(notplus[8]));
   INV_X1 i_1_9 (.A(secondVal[9]), .ZN(notplus[9]));
   INV_X1 i_1_10 (.A(secondVal[10]), .ZN(notplus[10]));
   INV_X1 i_1_11 (.A(secondVal[11]), .ZN(notplus[11]));
   INV_X1 i_1_12 (.A(secondVal[12]), .ZN(notplus[12]));
endmodule

module counterMux__22_29(counter, resetdata, dataIn, start, load, reset, 
      universalReset, continue, result);
   input [15:0]counter;
   input [15:0]resetdata;
   input [15:0]dataIn;
   input [15:0]start;
   input load;
   input reset;
   input universalReset;
   input continue;
   output [15:0]result;

   wire n_0_0;

   AND2_X1 i_0_0 (.A1(counter[0]), .A2(n_0_0), .ZN(result[0]));
   AND2_X1 i_0_1 (.A1(counter[1]), .A2(n_0_0), .ZN(result[1]));
   AND2_X1 i_0_2 (.A1(counter[2]), .A2(n_0_0), .ZN(result[2]));
   AND2_X1 i_0_3 (.A1(counter[3]), .A2(n_0_0), .ZN(result[3]));
   AND2_X1 i_0_4 (.A1(counter[4]), .A2(n_0_0), .ZN(result[4]));
   AND2_X1 i_0_5 (.A1(counter[5]), .A2(n_0_0), .ZN(result[5]));
   AND2_X1 i_0_6 (.A1(counter[6]), .A2(n_0_0), .ZN(result[6]));
   AND2_X1 i_0_7 (.A1(counter[7]), .A2(n_0_0), .ZN(result[7]));
   AND2_X1 i_0_8 (.A1(counter[8]), .A2(n_0_0), .ZN(result[8]));
   AND2_X1 i_0_9 (.A1(counter[9]), .A2(n_0_0), .ZN(result[9]));
   AND2_X1 i_0_10 (.A1(counter[10]), .A2(n_0_0), .ZN(result[10]));
   AND2_X1 i_0_11 (.A1(counter[11]), .A2(n_0_0), .ZN(result[11]));
   AND2_X1 i_0_12 (.A1(counter[12]), .A2(n_0_0), .ZN(result[12]));
   AND2_X1 i_0_13 (.A1(counter[13]), .A2(n_0_0), .ZN(result[13]));
   AND2_X1 i_0_14 (.A1(counter[14]), .A2(n_0_0), .ZN(result[14]));
   AND2_X1 i_0_15 (.A1(counter[15]), .A2(n_0_0), .ZN(result[15]));
   NOR2_X1 i_0_16 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
endmodule

module reg__22_26(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module counter__21_425(dataIn, offset, load, enable, CLK, reset, universalReset, 
      continue, dataOut, done, NFN);
   input [15:0]dataIn;
   input [15:0]offset;
   input load;
   input enable;
   input CLK;
   input reset;
   input universalReset;
   input continue;
   output [15:0]dataOut;
   output done;
   output NFN;

   wire [15:0]incremented;
   wire [15:0]muxOut;
   wire activate;
   wire n_0_0;
   wire n_0_1;

   Addition1__22_424 addition (.A(dataOut), .B(), .Cin(), .sum(incremented), 
      .overFlow());
   comparator__22_192 compare (.firstVal(dataOut), .secondVal({uc_0, uc_1, uc_2, 
      offset[12], offset[11], offset[10], offset[9], offset[8], offset[7], uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .done(n_0), .firstBigger(), 
      .firstSmaller());
   counterMux__22_29 muxing (.counter(incremented), .resetdata(), .dataIn(), 
      .start(), .load(), .reset(reset), .universalReset(universalReset), 
      .continue(), .result(muxOut));
   reg__22_26 count (.D(muxOut), .load(activate), .Clk(CLK), .Q(dataOut), 
      .rst(universalReset));
   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(n_0), .ZN(activate));
   NOR2_X1 i_0_1 (.A1(universalReset), .A2(reset), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(enable), .ZN(n_0_1));
endmodule

module mux__2_5005(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5008(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5011(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5014(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5017(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5020(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5023(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5026(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5029(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5032(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5035(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5038(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5041(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5044(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_0(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__2_2(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   mux__2_5005 muxx_1_muxx_j (.sel(B[0]), .in1(), .in2(), .i1(), .i2(B[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__2_5008 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(B[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__2_5011 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(B[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__2_5014 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(B[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__2_5017 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(B[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__2_5020 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(B[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__2_5023 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(B[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__2_5026 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(B[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__2_5029 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(B[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__2_5032 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(B[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__2_5035 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(B[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__2_5038 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(B[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__2_5041 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(B[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__2_5044 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(B[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__2_0 muxx_15_muxx_j (.sel(Carry), .in1(B[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module Partial_Full_Adder__2_601(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_597(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_593(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_589(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_585(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_581(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_577(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_573(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_569(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_565(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_561(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_557(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_553(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_549(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_545(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_541(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_634(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_601 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_597 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_593 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_589 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_585 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_581 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_577 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_573 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_569 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_565 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_561 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_557 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_553 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_549 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_545 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_541 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_769(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_765(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_761(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_757(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_753(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_749(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_745(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_741(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_737(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_733(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_729(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_725(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_721(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_717(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_713(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_709(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_802(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_769 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_765 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_761 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_757 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_753 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_749 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_745 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_741 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_737 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_733 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_729 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_725 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_721 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_717 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_713 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_709 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_937(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_933(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_929(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_925(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_921(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_917(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_913(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_909(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_905(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_901(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_897(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_893(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_889(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_885(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_881(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_877(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_970(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_937 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_933 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_929 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_925 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_921 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_917 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_913 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_909 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_905 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_901 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_897 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_893 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_889 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_885 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_881 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_877 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1105(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1101(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1097(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1093(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1089(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1085(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1081(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1077(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1073(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1069(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1065(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1061(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1057(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1053(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1049(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1045(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1138(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1105 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1101 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1097 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1093 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1089 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1085 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1081 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1077 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1073 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1069 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1065 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1061 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1057 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1053 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1049 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1045 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1273(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1269(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1265(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1261(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1257(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1253(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1249(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1245(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1241(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1237(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1233(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1229(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1225(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1221(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1217(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1213(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1306(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1273 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1269 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1265 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1261 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1257 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1253 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1249 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1245 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1241 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1237 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1233 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1229 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1225 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1221 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1217 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1213 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1441(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1437(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1433(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1429(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1425(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1421(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1417(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1413(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1409(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1405(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1401(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1397(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1393(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1389(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1385(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1381(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1474(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1441 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1437 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1433 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1429 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1425 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1421 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1417 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1413 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1409 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1405 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1401 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1397 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1393 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1389 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1385 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1381 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1609(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1605(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1601(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1597(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1593(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1589(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1585(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1581(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1577(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1573(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1569(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1565(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1561(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1557(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1553(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1549(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1642(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1609 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1605 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1601 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1597 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1593 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1589 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1585 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1581 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1577 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1573 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1569 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1565 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1561 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1557 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1553 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1549 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1777(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1773(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1769(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1765(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1761(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1757(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1753(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1749(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1745(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1741(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1737(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1733(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1729(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1725(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1721(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1717(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1810(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1777 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1773 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1769 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1765 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1761 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1757 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1753 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1749 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1745 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1741 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1737 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1733 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1729 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1725 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1721 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1717 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1945(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1941(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1937(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1933(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1929(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1925(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1921(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1917(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1913(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1909(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1905(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1901(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1897(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1893(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1889(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1885(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1978(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1945 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1941 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1937 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1933 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1929 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1925 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1921 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1917 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1913 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1909 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1905 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1901 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1897 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1893 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1889 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1885 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2113(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2109(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2105(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2101(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2097(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2093(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2089(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2085(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2081(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2077(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2073(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2069(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2065(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2061(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2057(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2053(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2146(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2113 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2109 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2105 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2101 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2097 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2093 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2089 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2085 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2081 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2077 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2073 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2069 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2065 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2061 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2057 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2053 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2281(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2277(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2273(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2269(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2265(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2261(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2257(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2253(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2249(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2245(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2241(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2237(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2233(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2229(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2225(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2221(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2314(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2281 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2277 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2273 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2269 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2265 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2261 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2257 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2253 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2249 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2245 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2241 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2237 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2233 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2229 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2225 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2221 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2449(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2445(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2441(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2437(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2433(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2429(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2425(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2421(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2417(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2413(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2409(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2405(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2401(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2397(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2393(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2389(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2482(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2449 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2445 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2441 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2437 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2433 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2429 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2425 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2421 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2417 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2413 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2409 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2405 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2401 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2397 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2393 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2389 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2617(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2613(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2609(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2605(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2601(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2597(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2593(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2589(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2585(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2581(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2577(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2573(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2569(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2565(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2561(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2557(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2650(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2617 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2613 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2609 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2605 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2601 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2597 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2593 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2589 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2585 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2581 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2577 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2573 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2569 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2565 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2561 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2557 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2785(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2781(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2777(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2773(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2769(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2765(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2761(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2757(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2753(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2749(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2745(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2741(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2737(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2733(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2729(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2725(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2818(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2785 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2781 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2777 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2773 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2769 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2765 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2761 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2757 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2753 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2749 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2745 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2741 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2737 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2733 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2729 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2725 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2953(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2949(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2945(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2941(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2937(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2933(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2929(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2925(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2921(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2917(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2913(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2909(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2905(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2901(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2897(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2893(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2986(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2953 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2949 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2945 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2941 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2937 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2933 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2929 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2925 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2921 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2917 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2913 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2909 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2905 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2901 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2897 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2893 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3121(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3117(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3113(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3109(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3105(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3101(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3097(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3093(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3089(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3085(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3081(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3077(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3073(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3069(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3065(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3061(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3154(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3121 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3117 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3113 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3109 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3105 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3101 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3097 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3093 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3089 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3085 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3081 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3077 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3073 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3069 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3065 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3061 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3289(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3285(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3281(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3277(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3273(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3269(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3265(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3261(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3257(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3253(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3249(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3245(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3241(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3237(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3233(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3229(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3322(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3289 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3285 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3281 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3277 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3273 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3269 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3265 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3261 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3257 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3253 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3249 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3245 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3241 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3237 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3233 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3229 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3457(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3453(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3449(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3445(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3441(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3437(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3433(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3429(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3425(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3421(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3417(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3413(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3409(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3405(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3401(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3397(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3490(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3457 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3453 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3449 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3445 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3441 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3437 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3433 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3429 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3425 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3421 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3417 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3413 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3409 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3405 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3401 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3397 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3625(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3621(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3617(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3613(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3609(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3605(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3601(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3597(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3593(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3589(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3585(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3581(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3577(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3573(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3569(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3565(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3658(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3625 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3621 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3617 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3613 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3609 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3605 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3601 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3597 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3593 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3589 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3585 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3581 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3577 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3573 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3569 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3565 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3793(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3789(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3785(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3781(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3777(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3773(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3769(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3765(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3761(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3757(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3753(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3749(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3745(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3741(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3737(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3733(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3826(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3793 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3789 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3785 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3781 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3777 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3773 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3769 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3765 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3761 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3757 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3753 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3749 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3745 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3741 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3737 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3733 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3961(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3957(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3953(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3949(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3945(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3941(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3937(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3933(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3929(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3925(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3921(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3917(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3913(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3909(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3905(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3901(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3994(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3961 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3957 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3953 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3949 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3945 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3941 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3937 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3933 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3929 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3925 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3921 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3917 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3913 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3909 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3905 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3901 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4129(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4125(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4121(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4117(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4113(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4109(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4105(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4101(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4097(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4093(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4089(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4085(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4081(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4077(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4073(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4069(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4162(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4129 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4125 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4121 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4117 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4113 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4109 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4105 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4101 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4097 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4093 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4089 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4085 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4081 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4077 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4073 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4069 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4297(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4293(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4289(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4285(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4281(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4277(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4273(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4269(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4265(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4261(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4257(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4253(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4249(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4245(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4241(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4237(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4330(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4297 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4293 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4289 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4285 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4281 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4277 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4273 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4269 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4265 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4261 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4257 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4253 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4249 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4245 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4241 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4237 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4465(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4461(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4457(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4453(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4449(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4445(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4441(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4437(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4433(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4429(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4425(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4421(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4417(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4413(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4409(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4405(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4498(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4465 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4461 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4457 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4453 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4449 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4445 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4441 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4437 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4433 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4429 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4425 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4421 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4417 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4413 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4409 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4405 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4633(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4629(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4625(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4621(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4617(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4613(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4609(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4605(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4601(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4597(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4593(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4589(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4585(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4581(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4577(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4573(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4666(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4633 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4629 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4625 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4621 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4617 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4613 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4609 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4605 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4601 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4597 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4593 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4589 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4585 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4581 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4577 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4573 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4801(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4797(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4793(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4789(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4785(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4781(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4777(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4773(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4769(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4765(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4761(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4757(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4753(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4749(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4745(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4741(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4834(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4801 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4797 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4793 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4789 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4785 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4781 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4777 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4773 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4769 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4765 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4761 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4757 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4753 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4749 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4745 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4741 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4969(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4965(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4961(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4957(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4953(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4949(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4945(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4941(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4937(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4933(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4929(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4925(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4921(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4917(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4913(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4909(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_5002(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_14;
   wire n_0_1;
   wire n_0_15;
   wire n_0_2;
   wire n_0_16;
   wire n_0_3;
   wire n_0_17;
   wire n_0_4;
   wire n_0_18;
   wire n_0_5;
   wire n_0_19;
   wire n_0_6;
   wire n_0_20;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4969 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4965 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_32), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4961 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_31), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4957 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_30), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4953 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_29), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4949 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_28), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4945 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_27), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4941 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(), .S(), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4937 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(), .S(), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4933 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(), .S(), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4929 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(), .S(), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4925 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(), .S(), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4921 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(), .S(), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4917 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(), .S(), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4913 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(), .S(), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4909 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_0_14));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_0_14), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_0_15));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_0_15), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_16));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_0_16), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_17));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_0_17), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_0_18));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_0_18), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_0_19));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_0_19), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_0_20));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_0_20), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_27));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_27), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_28));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_28), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_29));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_29), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_30));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_30), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_31));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_31), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_32));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_32), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_6(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_10(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_14(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_18(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_22(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_26(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_30(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_34(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_38(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_42(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_46(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_50(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_54(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_58(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_62(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_66(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_14;
   wire n_0_1;
   wire n_0_15;
   wire n_0_2;
   wire n_0_16;
   wire n_0_3;
   wire n_0_17;
   wire n_0_4;
   wire n_0_18;
   wire n_0_5;
   wire n_0_19;
   wire n_0_6;
   wire n_0_20;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_6 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_10 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_32), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_14 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_31), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_18 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_30), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_22 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_29), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_26 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_28), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_30 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_27), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_34 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(), .S(), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_38 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(), .S(), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_42 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(), .S(), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_46 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(), .S(), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_50 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(), .S(), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_54 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(), .S(), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_58 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(), .S(), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_62 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(), .S(), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_66 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_0_14));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_0_14), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_0_15));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_0_15), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_16));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_0_16), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_17));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_0_17), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_0_18));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_0_18), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_0_19));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_0_19), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_0_20));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_0_20), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_27));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_27), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_28));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_28), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_29));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_29), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_30));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_30), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_31));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_31), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_32));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_32), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module booth_multiplier(m, r, result, overflow);
   input [15:0]m;
   input [15:0]r;
   output [15:0]result;
   output overflow;

   wire [15:0]mn;
   wire [32:0]\temp1[1] ;
   wire [32:0]\temp2[1] ;
   wire [32:0]\temp1[2] ;
   wire [32:0]\temp2[2] ;
   wire [32:0]\temp1[3] ;
   wire [32:0]\temp2[3] ;
   wire [32:0]\temp1[4] ;
   wire [32:0]\temp2[4] ;
   wire [32:0]\temp1[5] ;
   wire [32:0]\temp2[5] ;
   wire [32:0]\temp1[6] ;
   wire [32:0]\temp2[6] ;
   wire [32:0]\temp1[7] ;
   wire [32:0]\temp2[7] ;
   wire [32:0]\temp1[8] ;
   wire [32:0]\temp2[8] ;
   wire [32:0]\temp1[9] ;
   wire [32:0]\temp2[9] ;
   wire [32:0]\temp1[10] ;
   wire [32:0]\temp2[10] ;
   wire [32:0]\temp1[11] ;
   wire [32:0]\temp2[11] ;
   wire [32:0]\temp1[12] ;
   wire [32:0]\temp2[12] ;
   wire [32:0]\temp1[13] ;
   wire [32:0]\temp2[13] ;
   wire [32:0]\temp2[14] ;
   wire [32:0]\temp1[14] ;
   wire [15:0]notM;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_177;
   wire n_1_178;
   wire n_1_179;
   wire n_1_180;
   wire n_1_181;
   wire n_1_182;
   wire n_1_183;
   wire n_1_184;
   wire n_1_185;
   wire n_1_186;
   wire n_1_187;
   wire n_1_188;
   wire n_1_189;
   wire n_1_190;
   wire n_1_191;
   wire n_1_192;
   wire n_1_193;
   wire n_1_194;
   wire n_1_195;
   wire n_1_196;
   wire n_1_197;
   wire n_1_198;
   wire n_1_199;
   wire n_1_200;
   wire n_1_201;
   wire n_1_202;
   wire n_1_203;
   wire n_1_204;
   wire n_1_205;
   wire n_1_206;
   wire n_1_207;
   wire n_1_208;
   wire n_1_209;
   wire n_1_210;
   wire n_1_211;
   wire n_1_212;
   wire n_1_213;
   wire n_1_214;
   wire n_1_215;
   wire n_1_216;
   wire n_1_217;
   wire n_1_218;
   wire n_1_219;
   wire n_1_220;
   wire n_1_221;
   wire n_1_222;
   wire n_1_223;
   wire n_1_224;
   wire n_1_225;
   wire n_1_226;
   wire n_1_227;
   wire n_1_228;
   wire n_1_229;
   wire n_1_230;
   wire n_1_231;
   wire n_1_232;
   wire n_1_233;
   wire n_1_234;
   wire n_1_235;
   wire n_1_236;
   wire n_1_237;
   wire n_1_238;
   wire n_1_239;
   wire n_1_240;
   wire n_1_241;
   wire n_1_242;
   wire n_1_243;
   wire n_1_244;
   wire n_1_245;
   wire n_1_246;
   wire n_1_247;
   wire n_1_248;
   wire n_1_249;
   wire n_1_250;
   wire n_1_251;
   wire n_1_252;
   wire n_1_253;
   wire n_1_254;
   wire n_1_255;
   wire n_1_256;
   wire n_1_257;
   wire n_1_258;
   wire n_1_259;
   wire n_1_260;
   wire n_1_261;
   wire n_1_262;
   wire n_1_263;
   wire n_1_264;
   wire n_1_265;
   wire n_1_266;
   wire n_1_267;
   wire n_1_268;
   wire n_1_269;
   wire n_1_270;
   wire n_1_271;
   wire n_1_272;
   wire n_1_273;
   wire n_1_274;
   wire n_1_275;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;

   Addition1__2_2 U0 (.A(), .B(notM), .Cin(), .sum({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], uc_0}), .overFlow());
   Carry_Look_Ahead_generic__2_634 x_1_Un (.A({n_209, uc_1, n_208, n_207, n_206, 
      n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, 
      n_195, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, 
      uc_13, uc_14, uc_15, uc_16, uc_17, uc_18}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, 
      uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35}), .Cin(), .S({
      \temp1[1] [32], \temp1[1] [31], \temp1[1] [30], \temp1[1] [29], 
      \temp1[1] [28], \temp1[1] [27], \temp1[1] [26], \temp1[1] [25], 
      \temp1[1] [24], \temp1[1] [23], \temp1[1] [22], \temp1[1] [21], 
      \temp1[1] [20], \temp1[1] [19], \temp1[1] [18], uc_36, uc_37, uc_38, uc_39, 
      uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, 
      uc_50, uc_51, uc_52, uc_53}), .overFlow());
   Carry_Look_Ahead_generic__2_802 x_1_Ux (.A({n_209, uc_54, n_208, n_207, n_206, 
      n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, 
      n_195, uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, 
      uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71}), .B({mn[15], 
      mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], 
      mn[4], mn[3], mn[2], mn[1], m[0], uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, 
      uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, 
      uc_88}), .Cin(), .S({\temp2[1] [32], \temp2[1] [31], \temp2[1] [30], 
      \temp2[1] [29], \temp2[1] [28], \temp2[1] [27], \temp2[1] [26], 
      \temp2[1] [25], \temp2[1] [24], \temp2[1] [23], \temp2[1] [22], 
      \temp2[1] [21], \temp2[1] [20], \temp2[1] [19], \temp2[1] [18], uc_89, 
      uc_90, uc_91, uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, uc_98, uc_99, 
      uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, uc_106}), .overFlow());
   Carry_Look_Ahead_generic__2_970 x_2_Un (.A({n_194, uc_107, n_193, n_192, 
      n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, 
      n_181, n_180, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, 
      uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, 
      uc_124}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_125, uc_126, uc_127, uc_128, 
      uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, 
      uc_138, uc_139, uc_140, uc_141}), .Cin(), .S({\temp1[2] [32], 
      \temp1[2] [31], \temp1[2] [30], \temp1[2] [29], \temp1[2] [28], 
      \temp1[2] [27], \temp1[2] [26], \temp1[2] [25], \temp1[2] [24], 
      \temp1[2] [23], \temp1[2] [22], \temp1[2] [21], \temp1[2] [20], 
      \temp1[2] [19], \temp1[2] [18], uc_142, uc_143, uc_144, uc_145, uc_146, 
      uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, uc_155, 
      uc_156, uc_157, uc_158, uc_159}), .overFlow());
   Carry_Look_Ahead_generic__2_1138 x_2_Ux (.A({n_194, uc_160, n_193, n_192, 
      n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, 
      n_181, n_180, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, 
      uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, 
      uc_177}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_178, uc_179, 
      uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, uc_186, uc_187, uc_188, 
      uc_189, uc_190, uc_191, uc_192, uc_193, uc_194}), .Cin(), .S({
      \temp2[2] [32], \temp2[2] [31], \temp2[2] [30], \temp2[2] [29], 
      \temp2[2] [28], \temp2[2] [27], \temp2[2] [26], \temp2[2] [25], 
      \temp2[2] [24], \temp2[2] [23], \temp2[2] [22], \temp2[2] [21], 
      \temp2[2] [20], \temp2[2] [19], \temp2[2] [18], uc_195, uc_196, uc_197, 
      uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, uc_204, uc_205, uc_206, 
      uc_207, uc_208, uc_209, uc_210, uc_211, uc_212}), .overFlow());
   Carry_Look_Ahead_generic__2_1306 x_3_Un (.A({n_179, uc_213, n_178, n_177, 
      n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
      n_166, n_165, uc_214, uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, 
      uc_221, uc_222, uc_223, uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, 
      uc_230}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_231, uc_232, uc_233, uc_234, 
      uc_235, uc_236, uc_237, uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, 
      uc_244, uc_245, uc_246, uc_247}), .Cin(), .S({\temp1[3] [32], 
      \temp1[3] [31], \temp1[3] [30], \temp1[3] [29], \temp1[3] [28], 
      \temp1[3] [27], \temp1[3] [26], \temp1[3] [25], \temp1[3] [24], 
      \temp1[3] [23], \temp1[3] [22], \temp1[3] [21], \temp1[3] [20], 
      \temp1[3] [19], \temp1[3] [18], uc_248, uc_249, uc_250, uc_251, uc_252, 
      uc_253, uc_254, uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, 
      uc_262, uc_263, uc_264, uc_265}), .overFlow());
   Carry_Look_Ahead_generic__2_1474 x_3_Ux (.A({n_179, uc_266, n_178, n_177, 
      n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
      n_166, n_165, uc_267, uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, 
      uc_274, uc_275, uc_276, uc_277, uc_278, uc_279, uc_280, uc_281, uc_282, 
      uc_283}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_284, uc_285, 
      uc_286, uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, uc_294, 
      uc_295, uc_296, uc_297, uc_298, uc_299, uc_300}), .Cin(), .S({
      \temp2[3] [32], \temp2[3] [31], \temp2[3] [30], \temp2[3] [29], 
      \temp2[3] [28], \temp2[3] [27], \temp2[3] [26], \temp2[3] [25], 
      \temp2[3] [24], \temp2[3] [23], \temp2[3] [22], \temp2[3] [21], 
      \temp2[3] [20], \temp2[3] [19], \temp2[3] [18], uc_301, uc_302, uc_303, 
      uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, 
      uc_313, uc_314, uc_315, uc_316, uc_317, uc_318}), .overFlow());
   Carry_Look_Ahead_generic__2_1642 x_4_Un (.A({n_164, uc_319, n_163, n_162, 
      n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, 
      n_151, n_150, uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, 
      uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, uc_334, uc_335, 
      uc_336}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_337, uc_338, uc_339, uc_340, 
      uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, uc_348, uc_349, 
      uc_350, uc_351, uc_352, uc_353}), .Cin(), .S({\temp1[4] [32], 
      \temp1[4] [31], \temp1[4] [30], \temp1[4] [29], \temp1[4] [28], 
      \temp1[4] [27], \temp1[4] [26], \temp1[4] [25], \temp1[4] [24], 
      \temp1[4] [23], \temp1[4] [22], \temp1[4] [21], \temp1[4] [20], 
      \temp1[4] [19], \temp1[4] [18], uc_354, uc_355, uc_356, uc_357, uc_358, 
      uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, uc_366, uc_367, 
      uc_368, uc_369, uc_370, uc_371}), .overFlow());
   Carry_Look_Ahead_generic__2_1810 x_4_Ux (.A({n_164, uc_372, n_163, n_162, 
      n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, 
      n_151, n_150, uc_373, uc_374, uc_375, uc_376, uc_377, uc_378, uc_379, 
      uc_380, uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, 
      uc_389}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_390, uc_391, 
      uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, uc_399, uc_400, 
      uc_401, uc_402, uc_403, uc_404, uc_405, uc_406}), .Cin(), .S({
      \temp2[4] [32], \temp2[4] [31], \temp2[4] [30], \temp2[4] [29], 
      \temp2[4] [28], \temp2[4] [27], \temp2[4] [26], \temp2[4] [25], 
      \temp2[4] [24], \temp2[4] [23], \temp2[4] [22], \temp2[4] [21], 
      \temp2[4] [20], \temp2[4] [19], \temp2[4] [18], uc_407, uc_408, uc_409, 
      uc_410, uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, 
      uc_419, uc_420, uc_421, uc_422, uc_423, uc_424}), .overFlow());
   Carry_Look_Ahead_generic__2_1978 x_5_Un (.A({n_149, uc_425, n_148, n_147, 
      n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
      n_136, n_135, uc_426, uc_427, uc_428, uc_429, uc_430, uc_431, uc_432, 
      uc_433, uc_434, uc_435, uc_436, uc_437, uc_438, uc_439, uc_440, uc_441, 
      uc_442}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_443, uc_444, uc_445, uc_446, 
      uc_447, uc_448, uc_449, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, 
      uc_456, uc_457, uc_458, uc_459}), .Cin(), .S({\temp1[5] [32], 
      \temp1[5] [31], \temp1[5] [30], \temp1[5] [29], \temp1[5] [28], 
      \temp1[5] [27], \temp1[5] [26], \temp1[5] [25], \temp1[5] [24], 
      \temp1[5] [23], \temp1[5] [22], \temp1[5] [21], \temp1[5] [20], 
      \temp1[5] [19], \temp1[5] [18], uc_460, uc_461, uc_462, uc_463, uc_464, 
      uc_465, uc_466, uc_467, uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, 
      uc_474, uc_475, uc_476, uc_477}), .overFlow());
   Carry_Look_Ahead_generic__2_2146 x_5_Ux (.A({n_149, uc_478, n_148, n_147, 
      n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
      n_136, n_135, uc_479, uc_480, uc_481, uc_482, uc_483, uc_484, uc_485, 
      uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, uc_492, uc_493, uc_494, 
      uc_495}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_496, uc_497, 
      uc_498, uc_499, uc_500, uc_501, uc_502, uc_503, uc_504, uc_505, uc_506, 
      uc_507, uc_508, uc_509, uc_510, uc_511, uc_512}), .Cin(), .S({
      \temp2[5] [32], \temp2[5] [31], \temp2[5] [30], \temp2[5] [29], 
      \temp2[5] [28], \temp2[5] [27], \temp2[5] [26], \temp2[5] [25], 
      \temp2[5] [24], \temp2[5] [23], \temp2[5] [22], \temp2[5] [21], 
      \temp2[5] [20], \temp2[5] [19], \temp2[5] [18], uc_513, uc_514, uc_515, 
      uc_516, uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, 
      uc_525, uc_526, uc_527, uc_528, uc_529, uc_530}), .overFlow());
   Carry_Look_Ahead_generic__2_2314 x_6_Un (.A({n_134, uc_531, n_133, n_132, 
      n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
      n_121, n_120, uc_532, uc_533, uc_534, uc_535, uc_536, uc_537, uc_538, 
      uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, uc_545, uc_546, uc_547, 
      uc_548}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_549, uc_550, uc_551, uc_552, 
      uc_553, uc_554, uc_555, uc_556, uc_557, uc_558, uc_559, uc_560, uc_561, 
      uc_562, uc_563, uc_564, uc_565}), .Cin(), .S({\temp1[6] [32], 
      \temp1[6] [31], \temp1[6] [30], \temp1[6] [29], \temp1[6] [28], 
      \temp1[6] [27], \temp1[6] [26], \temp1[6] [25], \temp1[6] [24], 
      \temp1[6] [23], \temp1[6] [22], \temp1[6] [21], \temp1[6] [20], 
      \temp1[6] [19], \temp1[6] [18], uc_566, uc_567, uc_568, uc_569, uc_570, 
      uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, 
      uc_580, uc_581, uc_582, uc_583}), .overFlow());
   Carry_Look_Ahead_generic__2_2482 x_6_Ux (.A({n_134, uc_584, n_133, n_132, 
      n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
      n_121, n_120, uc_585, uc_586, uc_587, uc_588, uc_589, uc_590, uc_591, 
      uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, uc_599, uc_600, 
      uc_601}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_602, uc_603, 
      uc_604, uc_605, uc_606, uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, 
      uc_613, uc_614, uc_615, uc_616, uc_617, uc_618}), .Cin(), .S({
      \temp2[6] [32], \temp2[6] [31], \temp2[6] [30], \temp2[6] [29], 
      \temp2[6] [28], \temp2[6] [27], \temp2[6] [26], \temp2[6] [25], 
      \temp2[6] [24], \temp2[6] [23], \temp2[6] [22], \temp2[6] [21], 
      \temp2[6] [20], \temp2[6] [19], \temp2[6] [18], uc_619, uc_620, uc_621, 
      uc_622, uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, uc_629, uc_630, 
      uc_631, uc_632, uc_633, uc_634, uc_635, uc_636}), .overFlow());
   Carry_Look_Ahead_generic__2_2650 x_7_Un (.A({n_119, uc_637, n_118, n_117, 
      n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
      n_106, n_105, uc_638, uc_639, uc_640, uc_641, uc_642, uc_643, uc_644, 
      uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, uc_651, uc_652, uc_653, 
      uc_654}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_655, uc_656, uc_657, uc_658, 
      uc_659, uc_660, uc_661, uc_662, uc_663, uc_664, uc_665, uc_666, uc_667, 
      uc_668, uc_669, uc_670, uc_671}), .Cin(), .S({\temp1[7] [32], 
      \temp1[7] [31], \temp1[7] [30], \temp1[7] [29], \temp1[7] [28], 
      \temp1[7] [27], \temp1[7] [26], \temp1[7] [25], \temp1[7] [24], 
      \temp1[7] [23], \temp1[7] [22], \temp1[7] [21], \temp1[7] [20], 
      \temp1[7] [19], \temp1[7] [18], uc_672, uc_673, uc_674, uc_675, uc_676, 
      uc_677, uc_678, uc_679, uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, 
      uc_686, uc_687, uc_688, uc_689}), .overFlow());
   Carry_Look_Ahead_generic__2_2818 x_7_Ux (.A({n_119, uc_690, n_118, n_117, 
      n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
      n_106, n_105, uc_691, uc_692, uc_693, uc_694, uc_695, uc_696, uc_697, 
      uc_698, uc_699, uc_700, uc_701, uc_702, uc_703, uc_704, uc_705, uc_706, 
      uc_707}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_708, uc_709, 
      uc_710, uc_711, uc_712, uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, 
      uc_719, uc_720, uc_721, uc_722, uc_723, uc_724}), .Cin(), .S({
      \temp2[7] [32], \temp2[7] [31], \temp2[7] [30], \temp2[7] [29], 
      \temp2[7] [28], \temp2[7] [27], \temp2[7] [26], \temp2[7] [25], 
      \temp2[7] [24], \temp2[7] [23], \temp2[7] [22], \temp2[7] [21], 
      \temp2[7] [20], \temp2[7] [19], \temp2[7] [18], uc_725, uc_726, uc_727, 
      uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, uc_734, uc_735, uc_736, 
      uc_737, uc_738, uc_739, uc_740, uc_741, uc_742}), .overFlow());
   Carry_Look_Ahead_generic__2_2986 x_8_Un (.A({n_104, uc_743, n_103, n_102, 
      n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
      uc_744, uc_745, uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, 
      uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, uc_760}), .B({
      m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_761, uc_762, uc_763, uc_764, uc_765, 
      uc_766, uc_767, uc_768, uc_769, uc_770, uc_771, uc_772, uc_773, uc_774, 
      uc_775, uc_776, uc_777}), .Cin(), .S({\temp1[8] [32], \temp1[8] [31], 
      \temp1[8] [30], \temp1[8] [29], \temp1[8] [28], \temp1[8] [27], 
      \temp1[8] [26], \temp1[8] [25], \temp1[8] [24], \temp1[8] [23], 
      \temp1[8] [22], \temp1[8] [21], \temp1[8] [20], \temp1[8] [19], 
      \temp1[8] [18], uc_778, uc_779, uc_780, uc_781, uc_782, uc_783, uc_784, 
      uc_785, uc_786, uc_787, uc_788, uc_789, uc_790, uc_791, uc_792, uc_793, 
      uc_794, uc_795}), .overFlow());
   Carry_Look_Ahead_generic__2_3154 x_8_Ux (.A({n_104, uc_796, n_103, n_102, 
      n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
      uc_797, uc_798, uc_799, uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, 
      uc_806, uc_807, uc_808, uc_809, uc_810, uc_811, uc_812, uc_813}), .B({
      mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], 
      mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_814, uc_815, uc_816, uc_817, 
      uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, uc_826, 
      uc_827, uc_828, uc_829, uc_830}), .Cin(), .S({\temp2[8] [32], 
      \temp2[8] [31], \temp2[8] [30], \temp2[8] [29], \temp2[8] [28], 
      \temp2[8] [27], \temp2[8] [26], \temp2[8] [25], \temp2[8] [24], 
      \temp2[8] [23], \temp2[8] [22], \temp2[8] [21], \temp2[8] [20], 
      \temp2[8] [19], \temp2[8] [18], uc_831, uc_832, uc_833, uc_834, uc_835, 
      uc_836, uc_837, uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, uc_844, 
      uc_845, uc_846, uc_847, uc_848}), .overFlow());
   Carry_Look_Ahead_generic__2_3322 x_9_Un (.A({n_89, uc_849, n_88, n_87, n_86, 
      n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, uc_850, 
      uc_851, uc_852, uc_853, uc_854, uc_855, uc_856, uc_857, uc_858, uc_859, 
      uc_860, uc_861, uc_862, uc_863, uc_864, uc_865, uc_866}), .B({m[15], m[14], 
      m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], 
      m[1], m[0], uc_867, uc_868, uc_869, uc_870, uc_871, uc_872, uc_873, uc_874, 
      uc_875, uc_876, uc_877, uc_878, uc_879, uc_880, uc_881, uc_882, uc_883}), 
      .Cin(), .S({\temp1[9] [32], \temp1[9] [31], \temp1[9] [30], \temp1[9] [29], 
      \temp1[9] [28], \temp1[9] [27], \temp1[9] [26], \temp1[9] [25], 
      \temp1[9] [24], \temp1[9] [23], \temp1[9] [22], \temp1[9] [21], 
      \temp1[9] [20], \temp1[9] [19], \temp1[9] [18], uc_884, uc_885, uc_886, 
      uc_887, uc_888, uc_889, uc_890, uc_891, uc_892, uc_893, uc_894, uc_895, 
      uc_896, uc_897, uc_898, uc_899, uc_900, uc_901}), .overFlow());
   Carry_Look_Ahead_generic__2_3490 x_9_Ux (.A({n_89, uc_902, n_88, n_87, n_86, 
      n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, uc_903, 
      uc_904, uc_905, uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, uc_912, 
      uc_913, uc_914, uc_915, uc_916, uc_917, uc_918, uc_919}), .B({mn[15], 
      mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], 
      mn[4], mn[3], mn[2], mn[1], m[0], uc_920, uc_921, uc_922, uc_923, uc_924, 
      uc_925, uc_926, uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, uc_933, 
      uc_934, uc_935, uc_936}), .Cin(), .S({\temp2[9] [32], \temp2[9] [31], 
      \temp2[9] [30], \temp2[9] [29], \temp2[9] [28], \temp2[9] [27], 
      \temp2[9] [26], \temp2[9] [25], \temp2[9] [24], \temp2[9] [23], 
      \temp2[9] [22], \temp2[9] [21], \temp2[9] [20], \temp2[9] [19], 
      \temp2[9] [18], uc_937, uc_938, uc_939, uc_940, uc_941, uc_942, uc_943, 
      uc_944, uc_945, uc_946, uc_947, uc_948, uc_949, uc_950, uc_951, uc_952, 
      uc_953, uc_954}), .overFlow());
   Carry_Look_Ahead_generic__2_3658 x_10_Un (.A({n_74, uc_955, n_73, n_72, n_71, 
      n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, uc_956, 
      uc_957, uc_958, uc_959, uc_960, uc_961, uc_962, uc_963, uc_964, uc_965, 
      uc_966, uc_967, uc_968, uc_969, uc_970, uc_971, uc_972}), .B({m[15], m[14], 
      m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], 
      m[1], m[0], uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, uc_979, uc_980, 
      uc_981, uc_982, uc_983, uc_984, uc_985, uc_986, uc_987, uc_988, uc_989}), 
      .Cin(), .S({\temp1[10] [32], \temp1[10] [31], \temp1[10] [30], 
      \temp1[10] [29], \temp1[10] [28], \temp1[10] [27], \temp1[10] [26], 
      \temp1[10] [25], \temp1[10] [24], \temp1[10] [23], \temp1[10] [22], 
      \temp1[10] [21], \temp1[10] [20], \temp1[10] [19], \temp1[10] [18], uc_990, 
      uc_991, uc_992, uc_993, uc_994, uc_995, uc_996, uc_997, uc_998, uc_999, 
      uc_1000, uc_1001, uc_1002, uc_1003, uc_1004, uc_1005, uc_1006, uc_1007}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_3826 x_10_Ux (.A({n_74, uc_1008, n_73, n_72, n_71, 
      n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, uc_1009, 
      uc_1010, uc_1011, uc_1012, uc_1013, uc_1014, uc_1015, uc_1016, uc_1017, 
      uc_1018, uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, uc_1024, uc_1025}), 
      .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], 
      mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1026, uc_1027, uc_1028, 
      uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, uc_1034, uc_1035, uc_1036, 
      uc_1037, uc_1038, uc_1039, uc_1040, uc_1041, uc_1042}), .Cin(), .S({
      \temp2[10] [32], \temp2[10] [31], \temp2[10] [30], \temp2[10] [29], 
      \temp2[10] [28], \temp2[10] [27], \temp2[10] [26], \temp2[10] [25], 
      \temp2[10] [24], \temp2[10] [23], \temp2[10] [22], \temp2[10] [21], 
      \temp2[10] [20], \temp2[10] [19], \temp2[10] [18], uc_1043, uc_1044, 
      uc_1045, uc_1046, uc_1047, uc_1048, uc_1049, uc_1050, uc_1051, uc_1052, 
      uc_1053, uc_1054, uc_1055, uc_1056, uc_1057, uc_1058, uc_1059, uc_1060}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_3994 x_11_Un (.A({n_59, uc_1061, n_58, n_57, n_56, 
      n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, uc_1062, 
      uc_1063, uc_1064, uc_1065, uc_1066, uc_1067, uc_1068, uc_1069, uc_1070, 
      uc_1071, uc_1072, uc_1073, uc_1074, uc_1075, uc_1076, uc_1077, uc_1078}), 
      .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_1079, uc_1080, uc_1081, uc_1082, uc_1083, 
      uc_1084, uc_1085, uc_1086, uc_1087, uc_1088, uc_1089, uc_1090, uc_1091, 
      uc_1092, uc_1093, uc_1094, uc_1095}), .Cin(), .S({\temp1[11] [32], 
      \temp1[11] [31], \temp1[11] [30], \temp1[11] [29], \temp1[11] [28], 
      \temp1[11] [27], \temp1[11] [26], \temp1[11] [25], \temp1[11] [24], 
      \temp1[11] [23], \temp1[11] [22], \temp1[11] [21], \temp1[11] [20], 
      \temp1[11] [19], \temp1[11] [18], uc_1096, uc_1097, uc_1098, uc_1099, 
      uc_1100, uc_1101, uc_1102, uc_1103, uc_1104, uc_1105, uc_1106, uc_1107, 
      uc_1108, uc_1109, uc_1110, uc_1111, uc_1112, uc_1113}), .overFlow());
   Carry_Look_Ahead_generic__2_4162 x_11_Ux (.A({n_59, uc_1114, n_58, n_57, n_56, 
      n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, uc_1115, 
      uc_1116, uc_1117, uc_1118, uc_1119, uc_1120, uc_1121, uc_1122, uc_1123, 
      uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, uc_1130, uc_1131}), 
      .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], 
      mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1132, uc_1133, uc_1134, 
      uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, uc_1140, uc_1141, uc_1142, 
      uc_1143, uc_1144, uc_1145, uc_1146, uc_1147, uc_1148}), .Cin(), .S({
      \temp2[11] [32], \temp2[11] [31], \temp2[11] [30], \temp2[11] [29], 
      \temp2[11] [28], \temp2[11] [27], \temp2[11] [26], \temp2[11] [25], 
      \temp2[11] [24], \temp2[11] [23], \temp2[11] [22], \temp2[11] [21], 
      \temp2[11] [20], \temp2[11] [19], \temp2[11] [18], uc_1149, uc_1150, 
      uc_1151, uc_1152, uc_1153, uc_1154, uc_1155, uc_1156, uc_1157, uc_1158, 
      uc_1159, uc_1160, uc_1161, uc_1162, uc_1163, uc_1164, uc_1165, uc_1166}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_4330 x_12_Un (.A({n_44, uc_1167, n_43, n_42, n_41, 
      n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, uc_1168, 
      uc_1169, uc_1170, uc_1171, uc_1172, uc_1173, uc_1174, uc_1175, uc_1176, 
      uc_1177, uc_1178, uc_1179, uc_1180, uc_1181, uc_1182, uc_1183, uc_1184}), 
      .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_1185, uc_1186, uc_1187, uc_1188, uc_1189, 
      uc_1190, uc_1191, uc_1192, uc_1193, uc_1194, uc_1195, uc_1196, uc_1197, 
      uc_1198, uc_1199, uc_1200, uc_1201}), .Cin(), .S({\temp1[12] [32], 
      \temp1[12] [31], \temp1[12] [30], \temp1[12] [29], \temp1[12] [28], 
      \temp1[12] [27], \temp1[12] [26], \temp1[12] [25], \temp1[12] [24], 
      \temp1[12] [23], \temp1[12] [22], \temp1[12] [21], \temp1[12] [20], 
      \temp1[12] [19], \temp1[12] [18], uc_1202, uc_1203, uc_1204, uc_1205, 
      uc_1206, uc_1207, uc_1208, uc_1209, uc_1210, uc_1211, uc_1212, uc_1213, 
      uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219}), .overFlow());
   Carry_Look_Ahead_generic__2_4498 x_12_Ux (.A({n_44, uc_1220, n_43, n_42, n_41, 
      n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, uc_1221, 
      uc_1222, uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, uc_1228, uc_1229, 
      uc_1230, uc_1231, uc_1232, uc_1233, uc_1234, uc_1235, uc_1236, uc_1237}), 
      .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], 
      mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1238, uc_1239, uc_1240, 
      uc_1241, uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, uc_1247, uc_1248, 
      uc_1249, uc_1250, uc_1251, uc_1252, uc_1253, uc_1254}), .Cin(), .S({
      \temp2[12] [32], \temp2[12] [31], \temp2[12] [30], \temp2[12] [29], 
      \temp2[12] [28], \temp2[12] [27], \temp2[12] [26], \temp2[12] [25], 
      \temp2[12] [24], \temp2[12] [23], \temp2[12] [22], \temp2[12] [21], 
      \temp2[12] [20], \temp2[12] [19], \temp2[12] [18], uc_1255, uc_1256, 
      uc_1257, uc_1258, uc_1259, uc_1260, uc_1261, uc_1262, uc_1263, uc_1264, 
      uc_1265, uc_1266, uc_1267, uc_1268, uc_1269, uc_1270, uc_1271, uc_1272}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_4666 x_13_Un (.A({n_29, uc_1273, n_28, n_27, n_26, 
      n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, uc_1274, 
      uc_1275, uc_1276, uc_1277, uc_1278, uc_1279, uc_1280, uc_1281, uc_1282, 
      uc_1283, uc_1284, uc_1285, uc_1286, uc_1287, uc_1288, uc_1289, uc_1290}), 
      .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_1291, uc_1292, uc_1293, uc_1294, uc_1295, 
      uc_1296, uc_1297, uc_1298, uc_1299, uc_1300, uc_1301, uc_1302, uc_1303, 
      uc_1304, uc_1305, uc_1306, uc_1307}), .Cin(), .S({\temp1[13] [32], 
      \temp1[13] [31], \temp1[13] [30], \temp1[13] [29], \temp1[13] [28], 
      \temp1[13] [27], \temp1[13] [26], \temp1[13] [25], \temp1[13] [24], 
      \temp1[13] [23], \temp1[13] [22], \temp1[13] [21], \temp1[13] [20], 
      \temp1[13] [19], \temp1[13] [18], uc_1308, uc_1309, uc_1310, uc_1311, 
      uc_1312, uc_1313, uc_1314, uc_1315, uc_1316, uc_1317, uc_1318, uc_1319, 
      uc_1320, uc_1321, uc_1322, uc_1323, uc_1324, uc_1325}), .overFlow());
   Carry_Look_Ahead_generic__2_4834 x_13_Ux (.A({n_29, uc_1326, n_28, n_27, n_26, 
      n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, uc_1327, 
      uc_1328, uc_1329, uc_1330, uc_1331, uc_1332, uc_1333, uc_1334, uc_1335, 
      uc_1336, uc_1337, uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, uc_1343}), 
      .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], 
      mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1344, uc_1345, uc_1346, 
      uc_1347, uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, uc_1353, uc_1354, 
      uc_1355, uc_1356, uc_1357, uc_1358, uc_1359, uc_1360}), .Cin(), .S({
      \temp2[13] [32], \temp2[13] [31], \temp2[13] [30], \temp2[13] [29], 
      \temp2[13] [28], \temp2[13] [27], \temp2[13] [26], \temp2[13] [25], 
      \temp2[13] [24], \temp2[13] [23], \temp2[13] [22], \temp2[13] [21], 
      \temp2[13] [20], \temp2[13] [19], \temp2[13] [18], uc_1361, uc_1362, 
      uc_1363, uc_1364, uc_1365, uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, 
      uc_1371, uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, uc_1378}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_5002 x_14_Ux (.A({n_14, uc_1379, n_13, n_12, n_11, 
      n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_1380, uc_1381, 
      uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, uc_1388, uc_1389, 
      uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396}), .B({
      mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], 
      mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1397, uc_1398, uc_1399, 
      uc_1400, uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, uc_1406, uc_1407, 
      uc_1408, uc_1409, uc_1410, uc_1411, uc_1412, uc_1413}), .Cin(), .S({
      \temp2[14] [32], \temp2[14] [31], \temp2[14] [30], \temp2[14] [29], 
      \temp2[14] [28], \temp2[14] [27], \temp2[14] [26], uc_1414, uc_1415, 
      uc_1416, uc_1417, uc_1418, uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, 
      uc_1424, uc_1425, uc_1426, uc_1427, uc_1428, uc_1429, uc_1430, uc_1431, 
      uc_1432, uc_1433, uc_1434, uc_1435, uc_1436, uc_1437, uc_1438, uc_1439}), 
      .overFlow());
   Carry_Look_Ahead_generic x_14_Un (.A({n_14, uc_1440, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_1441, uc_1442, 
      uc_1443, uc_1444, uc_1445, uc_1446, uc_1447, uc_1448, uc_1449, uc_1450, 
      uc_1451, uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, uc_1457}), .B({m[15], 
      m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], 
      m[3], m[2], m[1], m[0], uc_1458, uc_1459, uc_1460, uc_1461, uc_1462, 
      uc_1463, uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, uc_1469, uc_1470, 
      uc_1471, uc_1472, uc_1473, uc_1474}), .Cin(), .S({\temp1[14] [32], 
      \temp1[14] [31], \temp1[14] [30], \temp1[14] [29], \temp1[14] [28], 
      \temp1[14] [27], \temp1[14] [26], uc_1475, uc_1476, uc_1477, uc_1478, 
      uc_1479, uc_1480, uc_1481, uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, 
      uc_1487, uc_1488, uc_1489, uc_1490, uc_1491, uc_1492, uc_1493, uc_1494, 
      uc_1495, uc_1496, uc_1497, uc_1498, uc_1499, uc_1500}), .overFlow());
   INV_X1 i_0_0 (.A(m[0]), .ZN(notM[0]));
   INV_X1 i_0_1 (.A(m[1]), .ZN(notM[1]));
   INV_X1 i_0_2 (.A(m[2]), .ZN(notM[2]));
   INV_X1 i_0_3 (.A(m[3]), .ZN(notM[3]));
   INV_X1 i_0_4 (.A(m[4]), .ZN(notM[4]));
   INV_X1 i_0_5 (.A(m[5]), .ZN(notM[5]));
   INV_X1 i_0_6 (.A(m[6]), .ZN(notM[6]));
   INV_X1 i_0_7 (.A(m[7]), .ZN(notM[7]));
   INV_X1 i_0_8 (.A(m[8]), .ZN(notM[8]));
   INV_X1 i_0_9 (.A(m[9]), .ZN(notM[9]));
   INV_X1 i_0_10 (.A(m[10]), .ZN(notM[10]));
   INV_X1 i_0_11 (.A(m[11]), .ZN(notM[11]));
   INV_X1 i_0_12 (.A(m[12]), .ZN(notM[12]));
   INV_X1 i_0_13 (.A(m[13]), .ZN(notM[13]));
   INV_X1 i_0_14 (.A(m[14]), .ZN(notM[14]));
   INV_X1 i_0_15 (.A(m[15]), .ZN(notM[15]));
   AOI22_X1 i_1_0 (.A1(n_1_3), .A2(n_1_2), .B1(n_1_1), .B2(n_1_0), .ZN(overflow));
   NOR3_X1 i_1_1 (.A1(n_1_9), .A2(n_1_4), .A3(n_1_5), .ZN(n_1_0));
   NOR4_X1 i_1_2 (.A1(n_1_11), .A2(n_1_6), .A3(n_1_8), .A4(n_1_7), .ZN(n_1_1));
   AND3_X1 i_1_3 (.A1(n_1_9), .A2(n_1_7), .A3(n_1_6), .ZN(n_1_2));
   AND4_X1 i_1_4 (.A1(n_1_8), .A2(n_1_4), .A3(n_1_11), .A4(n_1_5), .ZN(n_1_3));
   AOI222_X1 i_1_5 (.A1(\temp1[14] [28]), .A2(n_1_30), .B1(\temp2[14] [28]), 
      .B2(n_1_29), .C1(n_11), .C2(n_1_28), .ZN(n_1_4));
   AOI222_X1 i_1_6 (.A1(\temp1[14] [27]), .A2(n_1_30), .B1(\temp2[14] [27]), 
      .B2(n_1_29), .C1(n_10), .C2(n_1_28), .ZN(n_1_5));
   AOI222_X1 i_1_7 (.A1(\temp1[14] [30]), .A2(n_1_30), .B1(\temp2[14] [30]), 
      .B2(n_1_29), .C1(n_13), .C2(n_1_28), .ZN(n_1_6));
   AOI222_X1 i_1_8 (.A1(\temp1[14] [29]), .A2(n_1_30), .B1(\temp2[14] [29]), 
      .B2(n_1_29), .C1(n_12), .C2(n_1_28), .ZN(n_1_7));
   AOI221_X1 i_1_9 (.A(n_1_10), .B1(\temp1[14] [31]), .B2(n_1_30), .C1(
      \temp2[14] [31]), .C2(n_1_29), .ZN(n_1_8));
   AOI221_X1 i_1_10 (.A(n_1_10), .B1(\temp1[14] [32]), .B2(n_1_30), .C1(
      \temp2[14] [32]), .C2(n_1_29), .ZN(n_1_9));
   AND2_X1 i_1_11 (.A1(n_14), .A2(n_1_28), .ZN(n_1_10));
   AOI222_X1 i_1_12 (.A1(\temp1[14] [26]), .A2(n_1_30), .B1(\temp2[14] [26]), 
      .B2(n_1_29), .C1(n_9), .C2(n_1_28), .ZN(n_1_11));
   NOR2_X1 i_1_45 (.A1(n_1_30), .A2(n_1_29), .ZN(n_1_28));
   AND2_X1 i_1_46 (.A1(r[14]), .A2(n_1_27), .ZN(n_1_29));
   NOR2_X1 i_1_47 (.A1(r[14]), .A2(n_1_27), .ZN(n_1_30));
   INV_X1 i_1_48 (.A(n_1_31), .ZN(n_0));
   AOI222_X1 i_1_49 (.A1(\temp1[13] [18]), .A2(n_1_49), .B1(\temp2[13] [18]), 
      .B2(n_1_48), .C1(n_16), .C2(n_1_47), .ZN(n_1_31));
   INV_X1 i_1_50 (.A(n_1_32), .ZN(n_1));
   AOI222_X1 i_1_51 (.A1(\temp1[13] [19]), .A2(n_1_49), .B1(\temp2[13] [19]), 
      .B2(n_1_48), .C1(n_17), .C2(n_1_47), .ZN(n_1_32));
   INV_X1 i_1_52 (.A(n_1_33), .ZN(n_2));
   AOI222_X1 i_1_53 (.A1(\temp1[13] [20]), .A2(n_1_49), .B1(\temp2[13] [20]), 
      .B2(n_1_48), .C1(n_18), .C2(n_1_47), .ZN(n_1_33));
   INV_X1 i_1_54 (.A(n_1_34), .ZN(n_3));
   AOI222_X1 i_1_55 (.A1(\temp1[13] [21]), .A2(n_1_49), .B1(\temp2[13] [21]), 
      .B2(n_1_48), .C1(n_19), .C2(n_1_47), .ZN(n_1_34));
   INV_X1 i_1_56 (.A(n_1_35), .ZN(n_4));
   AOI222_X1 i_1_57 (.A1(\temp1[13] [22]), .A2(n_1_49), .B1(\temp2[13] [22]), 
      .B2(n_1_48), .C1(n_20), .C2(n_1_47), .ZN(n_1_35));
   INV_X1 i_1_58 (.A(n_1_36), .ZN(n_5));
   AOI222_X1 i_1_59 (.A1(\temp1[13] [23]), .A2(n_1_49), .B1(\temp2[13] [23]), 
      .B2(n_1_48), .C1(n_21), .C2(n_1_47), .ZN(n_1_36));
   INV_X1 i_1_60 (.A(n_1_37), .ZN(n_6));
   AOI222_X1 i_1_61 (.A1(\temp1[13] [24]), .A2(n_1_49), .B1(\temp2[13] [24]), 
      .B2(n_1_48), .C1(n_22), .C2(n_1_47), .ZN(n_1_37));
   INV_X1 i_1_62 (.A(n_1_38), .ZN(n_7));
   AOI222_X1 i_1_63 (.A1(\temp1[13] [25]), .A2(n_1_49), .B1(\temp2[13] [25]), 
      .B2(n_1_48), .C1(n_23), .C2(n_1_47), .ZN(n_1_38));
   INV_X1 i_1_64 (.A(n_1_39), .ZN(n_8));
   AOI222_X1 i_1_65 (.A1(\temp1[13] [26]), .A2(n_1_49), .B1(\temp2[13] [26]), 
      .B2(n_1_48), .C1(n_24), .C2(n_1_47), .ZN(n_1_39));
   INV_X1 i_1_66 (.A(n_1_40), .ZN(n_9));
   AOI222_X1 i_1_67 (.A1(\temp1[13] [27]), .A2(n_1_49), .B1(\temp2[13] [27]), 
      .B2(n_1_48), .C1(n_25), .C2(n_1_47), .ZN(n_1_40));
   INV_X1 i_1_68 (.A(n_1_41), .ZN(n_10));
   AOI222_X1 i_1_69 (.A1(\temp1[13] [28]), .A2(n_1_49), .B1(\temp2[13] [28]), 
      .B2(n_1_48), .C1(n_26), .C2(n_1_47), .ZN(n_1_41));
   INV_X1 i_1_70 (.A(n_1_42), .ZN(n_11));
   AOI222_X1 i_1_71 (.A1(\temp1[13] [29]), .A2(n_1_49), .B1(\temp2[13] [29]), 
      .B2(n_1_48), .C1(n_27), .C2(n_1_47), .ZN(n_1_42));
   INV_X1 i_1_72 (.A(n_1_43), .ZN(n_12));
   AOI222_X1 i_1_73 (.A1(\temp1[13] [30]), .A2(n_1_49), .B1(\temp2[13] [30]), 
      .B2(n_1_48), .C1(n_28), .C2(n_1_47), .ZN(n_1_43));
   INV_X1 i_1_74 (.A(n_1_44), .ZN(n_13));
   AOI221_X1 i_1_75 (.A(n_1_46), .B1(\temp1[13] [31]), .B2(n_1_49), .C1(
      \temp2[13] [31]), .C2(n_1_48), .ZN(n_1_44));
   INV_X1 i_1_76 (.A(n_1_45), .ZN(n_14));
   AOI221_X1 i_1_77 (.A(n_1_46), .B1(\temp1[13] [32]), .B2(n_1_49), .C1(
      \temp2[13] [32]), .C2(n_1_48), .ZN(n_1_45));
   AND2_X1 i_1_78 (.A1(n_29), .A2(n_1_47), .ZN(n_1_46));
   NOR2_X1 i_1_79 (.A1(n_1_49), .A2(n_1_48), .ZN(n_1_47));
   NOR2_X1 i_1_80 (.A1(n_1_27), .A2(r[12]), .ZN(n_1_48));
   NOR2_X1 i_1_81 (.A1(r[13]), .A2(n_1_26), .ZN(n_1_49));
   INV_X1 i_1_82 (.A(n_1_50), .ZN(n_15));
   AOI222_X1 i_1_83 (.A1(\temp1[12] [18]), .A2(n_1_68), .B1(\temp2[12] [18]), 
      .B2(n_1_67), .C1(n_31), .C2(n_1_66), .ZN(n_1_50));
   INV_X1 i_1_84 (.A(n_1_51), .ZN(n_16));
   AOI222_X1 i_1_85 (.A1(\temp1[12] [19]), .A2(n_1_68), .B1(\temp2[12] [19]), 
      .B2(n_1_67), .C1(n_32), .C2(n_1_66), .ZN(n_1_51));
   INV_X1 i_1_86 (.A(n_1_52), .ZN(n_17));
   AOI222_X1 i_1_87 (.A1(\temp1[12] [20]), .A2(n_1_68), .B1(\temp2[12] [20]), 
      .B2(n_1_67), .C1(n_33), .C2(n_1_66), .ZN(n_1_52));
   INV_X1 i_1_88 (.A(n_1_53), .ZN(n_18));
   AOI222_X1 i_1_89 (.A1(\temp1[12] [21]), .A2(n_1_68), .B1(\temp2[12] [21]), 
      .B2(n_1_67), .C1(n_34), .C2(n_1_66), .ZN(n_1_53));
   INV_X1 i_1_90 (.A(n_1_54), .ZN(n_19));
   AOI222_X1 i_1_91 (.A1(\temp1[12] [22]), .A2(n_1_68), .B1(\temp2[12] [22]), 
      .B2(n_1_67), .C1(n_35), .C2(n_1_66), .ZN(n_1_54));
   INV_X1 i_1_92 (.A(n_1_55), .ZN(n_20));
   AOI222_X1 i_1_93 (.A1(\temp1[12] [23]), .A2(n_1_68), .B1(\temp2[12] [23]), 
      .B2(n_1_67), .C1(n_36), .C2(n_1_66), .ZN(n_1_55));
   INV_X1 i_1_94 (.A(n_1_56), .ZN(n_21));
   AOI222_X1 i_1_95 (.A1(\temp1[12] [24]), .A2(n_1_68), .B1(\temp2[12] [24]), 
      .B2(n_1_67), .C1(n_37), .C2(n_1_66), .ZN(n_1_56));
   INV_X1 i_1_96 (.A(n_1_57), .ZN(n_22));
   AOI222_X1 i_1_97 (.A1(\temp1[12] [25]), .A2(n_1_68), .B1(\temp2[12] [25]), 
      .B2(n_1_67), .C1(n_38), .C2(n_1_66), .ZN(n_1_57));
   INV_X1 i_1_98 (.A(n_1_58), .ZN(n_23));
   AOI222_X1 i_1_99 (.A1(\temp1[12] [26]), .A2(n_1_68), .B1(\temp2[12] [26]), 
      .B2(n_1_67), .C1(n_39), .C2(n_1_66), .ZN(n_1_58));
   INV_X1 i_1_100 (.A(n_1_59), .ZN(n_24));
   AOI222_X1 i_1_101 (.A1(\temp1[12] [27]), .A2(n_1_68), .B1(\temp2[12] [27]), 
      .B2(n_1_67), .C1(n_40), .C2(n_1_66), .ZN(n_1_59));
   INV_X1 i_1_102 (.A(n_1_60), .ZN(n_25));
   AOI222_X1 i_1_103 (.A1(\temp1[12] [28]), .A2(n_1_68), .B1(\temp2[12] [28]), 
      .B2(n_1_67), .C1(n_41), .C2(n_1_66), .ZN(n_1_60));
   INV_X1 i_1_104 (.A(n_1_61), .ZN(n_26));
   AOI222_X1 i_1_105 (.A1(\temp1[12] [29]), .A2(n_1_68), .B1(\temp2[12] [29]), 
      .B2(n_1_67), .C1(n_42), .C2(n_1_66), .ZN(n_1_61));
   INV_X1 i_1_106 (.A(n_1_62), .ZN(n_27));
   AOI222_X1 i_1_107 (.A1(\temp1[12] [30]), .A2(n_1_68), .B1(\temp2[12] [30]), 
      .B2(n_1_67), .C1(n_43), .C2(n_1_66), .ZN(n_1_62));
   INV_X1 i_1_108 (.A(n_1_63), .ZN(n_28));
   AOI221_X1 i_1_109 (.A(n_1_65), .B1(\temp1[12] [31]), .B2(n_1_68), .C1(
      \temp2[12] [31]), .C2(n_1_67), .ZN(n_1_63));
   INV_X1 i_1_110 (.A(n_1_64), .ZN(n_29));
   AOI221_X1 i_1_111 (.A(n_1_65), .B1(\temp1[12] [32]), .B2(n_1_68), .C1(
      \temp2[12] [32]), .C2(n_1_67), .ZN(n_1_64));
   AND2_X1 i_1_112 (.A1(n_44), .A2(n_1_66), .ZN(n_1_65));
   NOR2_X1 i_1_113 (.A1(n_1_68), .A2(n_1_67), .ZN(n_1_66));
   NOR2_X1 i_1_114 (.A1(n_1_26), .A2(r[11]), .ZN(n_1_67));
   NOR2_X1 i_1_115 (.A1(r[12]), .A2(n_1_25), .ZN(n_1_68));
   INV_X1 i_1_116 (.A(n_1_69), .ZN(n_30));
   AOI222_X1 i_1_117 (.A1(\temp1[11] [18]), .A2(n_1_87), .B1(\temp2[11] [18]), 
      .B2(n_1_86), .C1(n_46), .C2(n_1_85), .ZN(n_1_69));
   INV_X1 i_1_118 (.A(n_1_70), .ZN(n_31));
   AOI222_X1 i_1_119 (.A1(\temp1[11] [19]), .A2(n_1_87), .B1(\temp2[11] [19]), 
      .B2(n_1_86), .C1(n_47), .C2(n_1_85), .ZN(n_1_70));
   INV_X1 i_1_120 (.A(n_1_71), .ZN(n_32));
   AOI222_X1 i_1_121 (.A1(\temp1[11] [20]), .A2(n_1_87), .B1(\temp2[11] [20]), 
      .B2(n_1_86), .C1(n_48), .C2(n_1_85), .ZN(n_1_71));
   INV_X1 i_1_122 (.A(n_1_72), .ZN(n_33));
   AOI222_X1 i_1_123 (.A1(\temp1[11] [21]), .A2(n_1_87), .B1(\temp2[11] [21]), 
      .B2(n_1_86), .C1(n_49), .C2(n_1_85), .ZN(n_1_72));
   INV_X1 i_1_124 (.A(n_1_73), .ZN(n_34));
   AOI222_X1 i_1_125 (.A1(\temp1[11] [22]), .A2(n_1_87), .B1(\temp2[11] [22]), 
      .B2(n_1_86), .C1(n_50), .C2(n_1_85), .ZN(n_1_73));
   INV_X1 i_1_126 (.A(n_1_74), .ZN(n_35));
   AOI222_X1 i_1_127 (.A1(\temp1[11] [23]), .A2(n_1_87), .B1(\temp2[11] [23]), 
      .B2(n_1_86), .C1(n_51), .C2(n_1_85), .ZN(n_1_74));
   INV_X1 i_1_128 (.A(n_1_75), .ZN(n_36));
   AOI222_X1 i_1_129 (.A1(\temp1[11] [24]), .A2(n_1_87), .B1(\temp2[11] [24]), 
      .B2(n_1_86), .C1(n_52), .C2(n_1_85), .ZN(n_1_75));
   INV_X1 i_1_130 (.A(n_1_76), .ZN(n_37));
   AOI222_X1 i_1_131 (.A1(\temp1[11] [25]), .A2(n_1_87), .B1(\temp2[11] [25]), 
      .B2(n_1_86), .C1(n_53), .C2(n_1_85), .ZN(n_1_76));
   INV_X1 i_1_132 (.A(n_1_77), .ZN(n_38));
   AOI222_X1 i_1_133 (.A1(\temp1[11] [26]), .A2(n_1_87), .B1(\temp2[11] [26]), 
      .B2(n_1_86), .C1(n_54), .C2(n_1_85), .ZN(n_1_77));
   INV_X1 i_1_134 (.A(n_1_78), .ZN(n_39));
   AOI222_X1 i_1_135 (.A1(\temp1[11] [27]), .A2(n_1_87), .B1(\temp2[11] [27]), 
      .B2(n_1_86), .C1(n_55), .C2(n_1_85), .ZN(n_1_78));
   INV_X1 i_1_136 (.A(n_1_79), .ZN(n_40));
   AOI222_X1 i_1_137 (.A1(\temp2[11] [28]), .A2(n_1_86), .B1(\temp1[11] [28]), 
      .B2(n_1_87), .C1(n_56), .C2(n_1_85), .ZN(n_1_79));
   INV_X1 i_1_138 (.A(n_1_80), .ZN(n_41));
   AOI222_X1 i_1_139 (.A1(\temp1[11] [29]), .A2(n_1_87), .B1(\temp2[11] [29]), 
      .B2(n_1_86), .C1(n_57), .C2(n_1_85), .ZN(n_1_80));
   INV_X1 i_1_140 (.A(n_1_81), .ZN(n_42));
   AOI222_X1 i_1_141 (.A1(\temp1[11] [30]), .A2(n_1_87), .B1(\temp2[11] [30]), 
      .B2(n_1_86), .C1(n_58), .C2(n_1_85), .ZN(n_1_81));
   INV_X1 i_1_142 (.A(n_1_82), .ZN(n_43));
   AOI221_X1 i_1_143 (.A(n_1_84), .B1(\temp1[11] [31]), .B2(n_1_87), .C1(
      \temp2[11] [31]), .C2(n_1_86), .ZN(n_1_82));
   INV_X1 i_1_144 (.A(n_1_83), .ZN(n_44));
   AOI221_X1 i_1_145 (.A(n_1_84), .B1(\temp1[11] [32]), .B2(n_1_87), .C1(
      \temp2[11] [32]), .C2(n_1_86), .ZN(n_1_83));
   AND2_X1 i_1_146 (.A1(n_59), .A2(n_1_85), .ZN(n_1_84));
   NOR2_X1 i_1_147 (.A1(n_1_87), .A2(n_1_86), .ZN(n_1_85));
   NOR2_X1 i_1_148 (.A1(n_1_25), .A2(r[10]), .ZN(n_1_86));
   NOR2_X1 i_1_149 (.A1(r[11]), .A2(n_1_24), .ZN(n_1_87));
   INV_X1 i_1_150 (.A(n_1_88), .ZN(n_45));
   AOI222_X1 i_1_151 (.A1(\temp2[10] [18]), .A2(n_1_105), .B1(\temp1[10] [18]), 
      .B2(n_1_106), .C1(n_61), .C2(n_1_104), .ZN(n_1_88));
   INV_X1 i_1_152 (.A(n_1_89), .ZN(n_46));
   AOI222_X1 i_1_153 (.A1(\temp1[10] [19]), .A2(n_1_106), .B1(\temp2[10] [19]), 
      .B2(n_1_105), .C1(n_62), .C2(n_1_104), .ZN(n_1_89));
   INV_X1 i_1_154 (.A(n_1_90), .ZN(n_47));
   AOI222_X1 i_1_155 (.A1(\temp1[10] [20]), .A2(n_1_106), .B1(\temp2[10] [20]), 
      .B2(n_1_105), .C1(n_63), .C2(n_1_104), .ZN(n_1_90));
   INV_X1 i_1_156 (.A(n_1_91), .ZN(n_48));
   AOI222_X1 i_1_157 (.A1(\temp1[10] [21]), .A2(n_1_106), .B1(\temp2[10] [21]), 
      .B2(n_1_105), .C1(n_64), .C2(n_1_104), .ZN(n_1_91));
   INV_X1 i_1_158 (.A(n_1_92), .ZN(n_49));
   AOI222_X1 i_1_159 (.A1(\temp1[10] [22]), .A2(n_1_106), .B1(\temp2[10] [22]), 
      .B2(n_1_105), .C1(n_65), .C2(n_1_104), .ZN(n_1_92));
   INV_X1 i_1_160 (.A(n_1_93), .ZN(n_50));
   AOI222_X1 i_1_161 (.A1(\temp1[10] [23]), .A2(n_1_106), .B1(\temp2[10] [23]), 
      .B2(n_1_105), .C1(n_66), .C2(n_1_104), .ZN(n_1_93));
   INV_X1 i_1_162 (.A(n_1_94), .ZN(n_51));
   AOI222_X1 i_1_163 (.A1(\temp1[10] [24]), .A2(n_1_106), .B1(\temp2[10] [24]), 
      .B2(n_1_105), .C1(n_67), .C2(n_1_104), .ZN(n_1_94));
   INV_X1 i_1_164 (.A(n_1_95), .ZN(n_52));
   AOI222_X1 i_1_165 (.A1(\temp1[10] [25]), .A2(n_1_106), .B1(\temp2[10] [25]), 
      .B2(n_1_105), .C1(n_68), .C2(n_1_104), .ZN(n_1_95));
   INV_X1 i_1_166 (.A(n_1_96), .ZN(n_53));
   AOI222_X1 i_1_167 (.A1(\temp1[10] [26]), .A2(n_1_106), .B1(\temp2[10] [26]), 
      .B2(n_1_105), .C1(n_69), .C2(n_1_104), .ZN(n_1_96));
   INV_X1 i_1_168 (.A(n_1_97), .ZN(n_54));
   AOI222_X1 i_1_169 (.A1(\temp1[10] [27]), .A2(n_1_106), .B1(\temp2[10] [27]), 
      .B2(n_1_105), .C1(n_70), .C2(n_1_104), .ZN(n_1_97));
   INV_X1 i_1_170 (.A(n_1_98), .ZN(n_55));
   AOI222_X1 i_1_171 (.A1(\temp2[10] [28]), .A2(n_1_105), .B1(\temp1[10] [28]), 
      .B2(n_1_106), .C1(n_71), .C2(n_1_104), .ZN(n_1_98));
   INV_X1 i_1_172 (.A(n_1_99), .ZN(n_56));
   AOI222_X1 i_1_173 (.A1(\temp2[10] [29]), .A2(n_1_105), .B1(\temp1[10] [29]), 
      .B2(n_1_106), .C1(n_72), .C2(n_1_104), .ZN(n_1_99));
   INV_X1 i_1_174 (.A(n_1_100), .ZN(n_57));
   AOI222_X1 i_1_175 (.A1(\temp1[10] [30]), .A2(n_1_106), .B1(\temp2[10] [30]), 
      .B2(n_1_105), .C1(n_73), .C2(n_1_104), .ZN(n_1_100));
   INV_X1 i_1_176 (.A(n_1_101), .ZN(n_58));
   AOI221_X1 i_1_177 (.A(n_1_103), .B1(\temp1[10] [31]), .B2(n_1_106), .C1(
      \temp2[10] [31]), .C2(n_1_105), .ZN(n_1_101));
   INV_X1 i_1_178 (.A(n_1_102), .ZN(n_59));
   AOI221_X1 i_1_179 (.A(n_1_103), .B1(\temp1[10] [32]), .B2(n_1_106), .C1(
      \temp2[10] [32]), .C2(n_1_105), .ZN(n_1_102));
   AND2_X1 i_1_180 (.A1(n_74), .A2(n_1_104), .ZN(n_1_103));
   NOR2_X1 i_1_181 (.A1(n_1_106), .A2(n_1_105), .ZN(n_1_104));
   NOR2_X1 i_1_182 (.A1(n_1_24), .A2(r[9]), .ZN(n_1_105));
   NOR2_X1 i_1_183 (.A1(r[10]), .A2(n_1_23), .ZN(n_1_106));
   INV_X1 i_1_184 (.A(n_1_107), .ZN(n_60));
   AOI222_X1 i_1_185 (.A1(\temp2[9] [18]), .A2(n_1_124), .B1(\temp1[9] [18]), 
      .B2(n_1_125), .C1(n_76), .C2(n_1_123), .ZN(n_1_107));
   INV_X1 i_1_186 (.A(n_1_108), .ZN(n_61));
   AOI222_X1 i_1_187 (.A1(\temp2[9] [19]), .A2(n_1_124), .B1(\temp1[9] [19]), 
      .B2(n_1_125), .C1(n_77), .C2(n_1_123), .ZN(n_1_108));
   INV_X1 i_1_188 (.A(n_1_109), .ZN(n_62));
   AOI222_X1 i_1_189 (.A1(\temp2[9] [20]), .A2(n_1_124), .B1(\temp1[9] [20]), 
      .B2(n_1_125), .C1(n_78), .C2(n_1_123), .ZN(n_1_109));
   INV_X1 i_1_190 (.A(n_1_110), .ZN(n_63));
   AOI222_X1 i_1_191 (.A1(\temp1[9] [21]), .A2(n_1_125), .B1(\temp2[9] [21]), 
      .B2(n_1_124), .C1(n_79), .C2(n_1_123), .ZN(n_1_110));
   INV_X1 i_1_192 (.A(n_1_111), .ZN(n_64));
   AOI222_X1 i_1_193 (.A1(\temp1[9] [22]), .A2(n_1_125), .B1(\temp2[9] [22]), 
      .B2(n_1_124), .C1(n_80), .C2(n_1_123), .ZN(n_1_111));
   INV_X1 i_1_194 (.A(n_1_112), .ZN(n_65));
   AOI222_X1 i_1_195 (.A1(\temp1[9] [23]), .A2(n_1_125), .B1(\temp2[9] [23]), 
      .B2(n_1_124), .C1(n_81), .C2(n_1_123), .ZN(n_1_112));
   INV_X1 i_1_196 (.A(n_1_113), .ZN(n_66));
   AOI222_X1 i_1_197 (.A1(\temp1[9] [24]), .A2(n_1_125), .B1(\temp2[9] [24]), 
      .B2(n_1_124), .C1(n_82), .C2(n_1_123), .ZN(n_1_113));
   INV_X1 i_1_198 (.A(n_1_114), .ZN(n_67));
   AOI222_X1 i_1_199 (.A1(\temp1[9] [25]), .A2(n_1_125), .B1(\temp2[9] [25]), 
      .B2(n_1_124), .C1(n_83), .C2(n_1_123), .ZN(n_1_114));
   INV_X1 i_1_200 (.A(n_1_115), .ZN(n_68));
   AOI222_X1 i_1_201 (.A1(\temp1[9] [26]), .A2(n_1_125), .B1(\temp2[9] [26]), 
      .B2(n_1_124), .C1(n_84), .C2(n_1_123), .ZN(n_1_115));
   INV_X1 i_1_202 (.A(n_1_116), .ZN(n_69));
   AOI222_X1 i_1_203 (.A1(\temp1[9] [27]), .A2(n_1_125), .B1(\temp2[9] [27]), 
      .B2(n_1_124), .C1(n_85), .C2(n_1_123), .ZN(n_1_116));
   INV_X1 i_1_204 (.A(n_1_117), .ZN(n_70));
   AOI222_X1 i_1_205 (.A1(\temp2[9] [28]), .A2(n_1_124), .B1(\temp1[9] [28]), 
      .B2(n_1_125), .C1(n_86), .C2(n_1_123), .ZN(n_1_117));
   INV_X1 i_1_206 (.A(n_1_118), .ZN(n_71));
   AOI222_X1 i_1_207 (.A1(\temp2[9] [29]), .A2(n_1_124), .B1(\temp1[9] [29]), 
      .B2(n_1_125), .C1(n_87), .C2(n_1_123), .ZN(n_1_118));
   INV_X1 i_1_208 (.A(n_1_119), .ZN(n_72));
   AOI222_X1 i_1_209 (.A1(\temp2[9] [30]), .A2(n_1_124), .B1(\temp1[9] [30]), 
      .B2(n_1_125), .C1(n_88), .C2(n_1_123), .ZN(n_1_119));
   INV_X1 i_1_210 (.A(n_1_120), .ZN(n_73));
   AOI221_X1 i_1_211 (.A(n_1_122), .B1(\temp1[9] [31]), .B2(n_1_125), .C1(
      \temp2[9] [31]), .C2(n_1_124), .ZN(n_1_120));
   INV_X1 i_1_212 (.A(n_1_121), .ZN(n_74));
   AOI221_X1 i_1_213 (.A(n_1_122), .B1(\temp1[9] [32]), .B2(n_1_125), .C1(
      \temp2[9] [32]), .C2(n_1_124), .ZN(n_1_121));
   AND2_X1 i_1_214 (.A1(n_89), .A2(n_1_123), .ZN(n_1_122));
   NOR2_X1 i_1_215 (.A1(n_1_125), .A2(n_1_124), .ZN(n_1_123));
   NOR2_X1 i_1_216 (.A1(n_1_23), .A2(r[8]), .ZN(n_1_124));
   NOR2_X1 i_1_217 (.A1(r[9]), .A2(n_1_22), .ZN(n_1_125));
   INV_X1 i_1_218 (.A(n_1_126), .ZN(n_75));
   AOI222_X1 i_1_219 (.A1(\temp2[8] [18]), .A2(n_1_143), .B1(\temp1[8] [18]), 
      .B2(n_1_144), .C1(n_91), .C2(n_1_142), .ZN(n_1_126));
   INV_X1 i_1_220 (.A(n_1_127), .ZN(n_76));
   AOI222_X1 i_1_221 (.A1(\temp2[8] [19]), .A2(n_1_143), .B1(\temp1[8] [19]), 
      .B2(n_1_144), .C1(n_92), .C2(n_1_142), .ZN(n_1_127));
   INV_X1 i_1_222 (.A(n_1_128), .ZN(n_77));
   AOI222_X1 i_1_223 (.A1(\temp2[8] [20]), .A2(n_1_143), .B1(\temp1[8] [20]), 
      .B2(n_1_144), .C1(n_93), .C2(n_1_142), .ZN(n_1_128));
   INV_X1 i_1_224 (.A(n_1_129), .ZN(n_78));
   AOI222_X1 i_1_225 (.A1(\temp2[8] [21]), .A2(n_1_143), .B1(\temp1[8] [21]), 
      .B2(n_1_144), .C1(n_94), .C2(n_1_142), .ZN(n_1_129));
   INV_X1 i_1_226 (.A(n_1_130), .ZN(n_79));
   AOI222_X1 i_1_227 (.A1(\temp1[8] [22]), .A2(n_1_144), .B1(\temp2[8] [22]), 
      .B2(n_1_143), .C1(n_95), .C2(n_1_142), .ZN(n_1_130));
   INV_X1 i_1_228 (.A(n_1_131), .ZN(n_80));
   AOI222_X1 i_1_229 (.A1(\temp1[8] [23]), .A2(n_1_144), .B1(\temp2[8] [23]), 
      .B2(n_1_143), .C1(n_96), .C2(n_1_142), .ZN(n_1_131));
   INV_X1 i_1_230 (.A(n_1_132), .ZN(n_81));
   AOI222_X1 i_1_231 (.A1(\temp1[8] [24]), .A2(n_1_144), .B1(\temp2[8] [24]), 
      .B2(n_1_143), .C1(n_97), .C2(n_1_142), .ZN(n_1_132));
   INV_X1 i_1_232 (.A(n_1_133), .ZN(n_82));
   AOI222_X1 i_1_233 (.A1(\temp1[8] [25]), .A2(n_1_144), .B1(\temp2[8] [25]), 
      .B2(n_1_143), .C1(n_98), .C2(n_1_142), .ZN(n_1_133));
   INV_X1 i_1_234 (.A(n_1_134), .ZN(n_83));
   AOI222_X1 i_1_235 (.A1(\temp1[8] [26]), .A2(n_1_144), .B1(\temp2[8] [26]), 
      .B2(n_1_143), .C1(n_99), .C2(n_1_142), .ZN(n_1_134));
   INV_X1 i_1_236 (.A(n_1_135), .ZN(n_84));
   AOI222_X1 i_1_237 (.A1(\temp1[8] [27]), .A2(n_1_144), .B1(\temp2[8] [27]), 
      .B2(n_1_143), .C1(n_100), .C2(n_1_142), .ZN(n_1_135));
   INV_X1 i_1_238 (.A(n_1_136), .ZN(n_85));
   AOI222_X1 i_1_239 (.A1(\temp2[8] [28]), .A2(n_1_143), .B1(\temp1[8] [28]), 
      .B2(n_1_144), .C1(n_101), .C2(n_1_142), .ZN(n_1_136));
   INV_X1 i_1_240 (.A(n_1_137), .ZN(n_86));
   AOI222_X1 i_1_241 (.A1(\temp2[8] [29]), .A2(n_1_143), .B1(\temp1[8] [29]), 
      .B2(n_1_144), .C1(n_102), .C2(n_1_142), .ZN(n_1_137));
   INV_X1 i_1_242 (.A(n_1_138), .ZN(n_87));
   AOI222_X1 i_1_243 (.A1(\temp2[8] [30]), .A2(n_1_143), .B1(\temp1[8] [30]), 
      .B2(n_1_144), .C1(n_103), .C2(n_1_142), .ZN(n_1_138));
   INV_X1 i_1_244 (.A(n_1_139), .ZN(n_88));
   AOI221_X1 i_1_245 (.A(n_1_141), .B1(\temp1[8] [31]), .B2(n_1_144), .C1(
      \temp2[8] [31]), .C2(n_1_143), .ZN(n_1_139));
   INV_X1 i_1_246 (.A(n_1_140), .ZN(n_89));
   AOI221_X1 i_1_247 (.A(n_1_141), .B1(\temp1[8] [32]), .B2(n_1_144), .C1(
      \temp2[8] [32]), .C2(n_1_143), .ZN(n_1_140));
   AND2_X1 i_1_248 (.A1(n_104), .A2(n_1_142), .ZN(n_1_141));
   NOR2_X1 i_1_249 (.A1(n_1_144), .A2(n_1_143), .ZN(n_1_142));
   NOR2_X1 i_1_250 (.A1(n_1_22), .A2(r[7]), .ZN(n_1_143));
   NOR2_X1 i_1_251 (.A1(r[8]), .A2(n_1_21), .ZN(n_1_144));
   INV_X1 i_1_252 (.A(n_1_145), .ZN(n_90));
   AOI222_X1 i_1_253 (.A1(\temp2[7] [18]), .A2(n_1_162), .B1(\temp1[7] [18]), 
      .B2(n_1_163), .C1(n_106), .C2(n_1_161), .ZN(n_1_145));
   INV_X1 i_1_254 (.A(n_1_146), .ZN(n_91));
   AOI222_X1 i_1_255 (.A1(\temp2[7] [19]), .A2(n_1_162), .B1(\temp1[7] [19]), 
      .B2(n_1_163), .C1(n_107), .C2(n_1_161), .ZN(n_1_146));
   INV_X1 i_1_256 (.A(n_1_147), .ZN(n_92));
   AOI222_X1 i_1_257 (.A1(\temp2[7] [20]), .A2(n_1_162), .B1(\temp1[7] [20]), 
      .B2(n_1_163), .C1(n_108), .C2(n_1_161), .ZN(n_1_147));
   INV_X1 i_1_258 (.A(n_1_148), .ZN(n_93));
   AOI222_X1 i_1_259 (.A1(\temp2[7] [21]), .A2(n_1_162), .B1(\temp1[7] [21]), 
      .B2(n_1_163), .C1(n_109), .C2(n_1_161), .ZN(n_1_148));
   INV_X1 i_1_260 (.A(n_1_149), .ZN(n_94));
   AOI222_X1 i_1_261 (.A1(\temp2[7] [22]), .A2(n_1_162), .B1(\temp1[7] [22]), 
      .B2(n_1_163), .C1(n_110), .C2(n_1_161), .ZN(n_1_149));
   INV_X1 i_1_262 (.A(n_1_150), .ZN(n_95));
   AOI222_X1 i_1_263 (.A1(\temp2[7] [23]), .A2(n_1_162), .B1(\temp1[7] [23]), 
      .B2(n_1_163), .C1(n_111), .C2(n_1_161), .ZN(n_1_150));
   INV_X1 i_1_264 (.A(n_1_151), .ZN(n_96));
   AOI222_X1 i_1_265 (.A1(\temp1[7] [24]), .A2(n_1_163), .B1(\temp2[7] [24]), 
      .B2(n_1_162), .C1(n_112), .C2(n_1_161), .ZN(n_1_151));
   INV_X1 i_1_266 (.A(n_1_152), .ZN(n_97));
   AOI222_X1 i_1_267 (.A1(\temp1[7] [25]), .A2(n_1_163), .B1(\temp2[7] [25]), 
      .B2(n_1_162), .C1(n_113), .C2(n_1_161), .ZN(n_1_152));
   INV_X1 i_1_268 (.A(n_1_153), .ZN(n_98));
   AOI222_X1 i_1_269 (.A1(\temp1[7] [26]), .A2(n_1_163), .B1(\temp2[7] [26]), 
      .B2(n_1_162), .C1(n_114), .C2(n_1_161), .ZN(n_1_153));
   INV_X1 i_1_270 (.A(n_1_154), .ZN(n_99));
   AOI222_X1 i_1_271 (.A1(\temp1[7] [27]), .A2(n_1_163), .B1(\temp2[7] [27]), 
      .B2(n_1_162), .C1(n_115), .C2(n_1_161), .ZN(n_1_154));
   INV_X1 i_1_272 (.A(n_1_155), .ZN(n_100));
   AOI222_X1 i_1_273 (.A1(\temp2[7] [28]), .A2(n_1_162), .B1(\temp1[7] [28]), 
      .B2(n_1_163), .C1(n_116), .C2(n_1_161), .ZN(n_1_155));
   INV_X1 i_1_274 (.A(n_1_156), .ZN(n_101));
   AOI222_X1 i_1_275 (.A1(\temp2[7] [29]), .A2(n_1_162), .B1(\temp1[7] [29]), 
      .B2(n_1_163), .C1(n_117), .C2(n_1_161), .ZN(n_1_156));
   INV_X1 i_1_276 (.A(n_1_157), .ZN(n_102));
   AOI222_X1 i_1_277 (.A1(\temp2[7] [30]), .A2(n_1_162), .B1(\temp1[7] [30]), 
      .B2(n_1_163), .C1(n_118), .C2(n_1_161), .ZN(n_1_157));
   INV_X1 i_1_278 (.A(n_1_158), .ZN(n_103));
   AOI221_X1 i_1_279 (.A(n_1_160), .B1(\temp1[7] [31]), .B2(n_1_163), .C1(
      \temp2[7] [31]), .C2(n_1_162), .ZN(n_1_158));
   INV_X1 i_1_280 (.A(n_1_159), .ZN(n_104));
   AOI221_X1 i_1_281 (.A(n_1_160), .B1(\temp1[7] [32]), .B2(n_1_163), .C1(
      \temp2[7] [32]), .C2(n_1_162), .ZN(n_1_159));
   AND2_X1 i_1_282 (.A1(n_119), .A2(n_1_161), .ZN(n_1_160));
   NOR2_X1 i_1_283 (.A1(n_1_163), .A2(n_1_162), .ZN(n_1_161));
   NOR2_X1 i_1_284 (.A1(n_1_21), .A2(r[6]), .ZN(n_1_162));
   NOR2_X1 i_1_285 (.A1(r[7]), .A2(n_1_20), .ZN(n_1_163));
   INV_X1 i_1_286 (.A(n_1_164), .ZN(n_105));
   AOI222_X1 i_1_287 (.A1(\temp2[6] [18]), .A2(n_1_181), .B1(\temp1[6] [18]), 
      .B2(n_1_182), .C1(n_121), .C2(n_1_180), .ZN(n_1_164));
   INV_X1 i_1_288 (.A(n_1_165), .ZN(n_106));
   AOI222_X1 i_1_289 (.A1(\temp2[6] [19]), .A2(n_1_181), .B1(\temp1[6] [19]), 
      .B2(n_1_182), .C1(n_122), .C2(n_1_180), .ZN(n_1_165));
   INV_X1 i_1_290 (.A(n_1_166), .ZN(n_107));
   AOI222_X1 i_1_291 (.A1(\temp2[6] [20]), .A2(n_1_181), .B1(\temp1[6] [20]), 
      .B2(n_1_182), .C1(n_123), .C2(n_1_180), .ZN(n_1_166));
   INV_X1 i_1_292 (.A(n_1_167), .ZN(n_108));
   AOI222_X1 i_1_293 (.A1(\temp2[6] [21]), .A2(n_1_181), .B1(\temp1[6] [21]), 
      .B2(n_1_182), .C1(n_124), .C2(n_1_180), .ZN(n_1_167));
   INV_X1 i_1_294 (.A(n_1_168), .ZN(n_109));
   AOI222_X1 i_1_295 (.A1(\temp2[6] [22]), .A2(n_1_181), .B1(\temp1[6] [22]), 
      .B2(n_1_182), .C1(n_125), .C2(n_1_180), .ZN(n_1_168));
   INV_X1 i_1_296 (.A(n_1_169), .ZN(n_110));
   AOI222_X1 i_1_297 (.A1(\temp2[6] [23]), .A2(n_1_181), .B1(\temp1[6] [23]), 
      .B2(n_1_182), .C1(n_126), .C2(n_1_180), .ZN(n_1_169));
   INV_X1 i_1_298 (.A(n_1_170), .ZN(n_111));
   AOI222_X1 i_1_299 (.A1(\temp2[6] [24]), .A2(n_1_181), .B1(\temp1[6] [24]), 
      .B2(n_1_182), .C1(n_127), .C2(n_1_180), .ZN(n_1_170));
   INV_X1 i_1_300 (.A(n_1_171), .ZN(n_112));
   AOI222_X1 i_1_301 (.A1(\temp1[6] [25]), .A2(n_1_182), .B1(\temp2[6] [25]), 
      .B2(n_1_181), .C1(n_128), .C2(n_1_180), .ZN(n_1_171));
   INV_X1 i_1_302 (.A(n_1_172), .ZN(n_113));
   AOI222_X1 i_1_303 (.A1(\temp1[6] [26]), .A2(n_1_182), .B1(\temp2[6] [26]), 
      .B2(n_1_181), .C1(n_129), .C2(n_1_180), .ZN(n_1_172));
   INV_X1 i_1_304 (.A(n_1_173), .ZN(n_114));
   AOI222_X1 i_1_305 (.A1(\temp1[6] [27]), .A2(n_1_182), .B1(\temp2[6] [27]), 
      .B2(n_1_181), .C1(n_130), .C2(n_1_180), .ZN(n_1_173));
   INV_X1 i_1_306 (.A(n_1_174), .ZN(n_115));
   AOI222_X1 i_1_307 (.A1(\temp2[6] [28]), .A2(n_1_181), .B1(\temp1[6] [28]), 
      .B2(n_1_182), .C1(n_131), .C2(n_1_180), .ZN(n_1_174));
   INV_X1 i_1_308 (.A(n_1_175), .ZN(n_116));
   AOI222_X1 i_1_309 (.A1(\temp2[6] [29]), .A2(n_1_181), .B1(\temp1[6] [29]), 
      .B2(n_1_182), .C1(n_132), .C2(n_1_180), .ZN(n_1_175));
   INV_X1 i_1_310 (.A(n_1_176), .ZN(n_117));
   AOI222_X1 i_1_311 (.A1(\temp2[6] [30]), .A2(n_1_181), .B1(\temp1[6] [30]), 
      .B2(n_1_182), .C1(n_133), .C2(n_1_180), .ZN(n_1_176));
   INV_X1 i_1_312 (.A(n_1_177), .ZN(n_118));
   AOI221_X1 i_1_313 (.A(n_1_179), .B1(\temp1[6] [31]), .B2(n_1_182), .C1(
      \temp2[6] [31]), .C2(n_1_181), .ZN(n_1_177));
   INV_X1 i_1_314 (.A(n_1_178), .ZN(n_119));
   AOI221_X1 i_1_315 (.A(n_1_179), .B1(\temp1[6] [32]), .B2(n_1_182), .C1(
      \temp2[6] [32]), .C2(n_1_181), .ZN(n_1_178));
   AND2_X1 i_1_316 (.A1(n_134), .A2(n_1_180), .ZN(n_1_179));
   NOR2_X1 i_1_317 (.A1(n_1_182), .A2(n_1_181), .ZN(n_1_180));
   NOR2_X1 i_1_318 (.A1(n_1_20), .A2(r[5]), .ZN(n_1_181));
   NOR2_X1 i_1_319 (.A1(r[6]), .A2(n_1_19), .ZN(n_1_182));
   INV_X1 i_1_320 (.A(n_1_183), .ZN(n_120));
   AOI222_X1 i_1_321 (.A1(\temp2[5] [18]), .A2(n_1_200), .B1(\temp1[5] [18]), 
      .B2(n_1_201), .C1(n_136), .C2(n_1_199), .ZN(n_1_183));
   INV_X1 i_1_322 (.A(n_1_184), .ZN(n_121));
   AOI222_X1 i_1_323 (.A1(\temp2[5] [19]), .A2(n_1_200), .B1(\temp1[5] [19]), 
      .B2(n_1_201), .C1(n_137), .C2(n_1_199), .ZN(n_1_184));
   INV_X1 i_1_324 (.A(n_1_185), .ZN(n_122));
   AOI222_X1 i_1_325 (.A1(\temp2[5] [20]), .A2(n_1_200), .B1(\temp1[5] [20]), 
      .B2(n_1_201), .C1(n_138), .C2(n_1_199), .ZN(n_1_185));
   INV_X1 i_1_326 (.A(n_1_186), .ZN(n_123));
   AOI222_X1 i_1_327 (.A1(\temp2[5] [21]), .A2(n_1_200), .B1(\temp1[5] [21]), 
      .B2(n_1_201), .C1(n_139), .C2(n_1_199), .ZN(n_1_186));
   INV_X1 i_1_328 (.A(n_1_187), .ZN(n_124));
   AOI222_X1 i_1_329 (.A1(\temp2[5] [22]), .A2(n_1_200), .B1(\temp1[5] [22]), 
      .B2(n_1_201), .C1(n_140), .C2(n_1_199), .ZN(n_1_187));
   INV_X1 i_1_330 (.A(n_1_188), .ZN(n_125));
   AOI222_X1 i_1_331 (.A1(\temp2[5] [23]), .A2(n_1_200), .B1(\temp1[5] [23]), 
      .B2(n_1_201), .C1(n_141), .C2(n_1_199), .ZN(n_1_188));
   INV_X1 i_1_332 (.A(n_1_189), .ZN(n_126));
   AOI222_X1 i_1_333 (.A1(\temp2[5] [24]), .A2(n_1_200), .B1(\temp1[5] [24]), 
      .B2(n_1_201), .C1(n_142), .C2(n_1_199), .ZN(n_1_189));
   INV_X1 i_1_334 (.A(n_1_190), .ZN(n_127));
   AOI222_X1 i_1_335 (.A1(\temp2[5] [25]), .A2(n_1_200), .B1(\temp1[5] [25]), 
      .B2(n_1_201), .C1(n_143), .C2(n_1_199), .ZN(n_1_190));
   INV_X1 i_1_336 (.A(n_1_191), .ZN(n_128));
   AOI222_X1 i_1_337 (.A1(\temp2[5] [26]), .A2(n_1_200), .B1(\temp1[5] [26]), 
      .B2(n_1_201), .C1(n_144), .C2(n_1_199), .ZN(n_1_191));
   INV_X1 i_1_338 (.A(n_1_192), .ZN(n_129));
   AOI222_X1 i_1_339 (.A1(\temp2[5] [27]), .A2(n_1_200), .B1(\temp1[5] [27]), 
      .B2(n_1_201), .C1(n_145), .C2(n_1_199), .ZN(n_1_192));
   INV_X1 i_1_340 (.A(n_1_193), .ZN(n_130));
   AOI222_X1 i_1_341 (.A1(\temp2[5] [28]), .A2(n_1_200), .B1(\temp1[5] [28]), 
      .B2(n_1_201), .C1(n_146), .C2(n_1_199), .ZN(n_1_193));
   INV_X1 i_1_342 (.A(n_1_194), .ZN(n_131));
   AOI222_X1 i_1_343 (.A1(\temp2[5] [29]), .A2(n_1_200), .B1(\temp1[5] [29]), 
      .B2(n_1_201), .C1(n_147), .C2(n_1_199), .ZN(n_1_194));
   INV_X1 i_1_344 (.A(n_1_195), .ZN(n_132));
   AOI222_X1 i_1_345 (.A1(\temp2[5] [30]), .A2(n_1_200), .B1(\temp1[5] [30]), 
      .B2(n_1_201), .C1(n_148), .C2(n_1_199), .ZN(n_1_195));
   INV_X1 i_1_346 (.A(n_1_196), .ZN(n_133));
   AOI221_X1 i_1_347 (.A(n_1_198), .B1(\temp1[5] [31]), .B2(n_1_201), .C1(
      \temp2[5] [31]), .C2(n_1_200), .ZN(n_1_196));
   INV_X1 i_1_348 (.A(n_1_197), .ZN(n_134));
   AOI221_X1 i_1_349 (.A(n_1_198), .B1(\temp1[5] [32]), .B2(n_1_201), .C1(
      \temp2[5] [32]), .C2(n_1_200), .ZN(n_1_197));
   AND2_X1 i_1_350 (.A1(n_149), .A2(n_1_199), .ZN(n_1_198));
   NOR2_X1 i_1_351 (.A1(n_1_201), .A2(n_1_200), .ZN(n_1_199));
   NOR2_X1 i_1_352 (.A1(n_1_19), .A2(r[4]), .ZN(n_1_200));
   NOR2_X1 i_1_353 (.A1(r[5]), .A2(n_1_18), .ZN(n_1_201));
   INV_X1 i_1_354 (.A(n_1_202), .ZN(n_135));
   AOI222_X1 i_1_355 (.A1(\temp2[4] [18]), .A2(n_1_219), .B1(\temp1[4] [18]), 
      .B2(n_1_220), .C1(n_151), .C2(n_1_218), .ZN(n_1_202));
   INV_X1 i_1_356 (.A(n_1_203), .ZN(n_136));
   AOI222_X1 i_1_357 (.A1(\temp2[4] [19]), .A2(n_1_219), .B1(\temp1[4] [19]), 
      .B2(n_1_220), .C1(n_152), .C2(n_1_218), .ZN(n_1_203));
   INV_X1 i_1_358 (.A(n_1_204), .ZN(n_137));
   AOI222_X1 i_1_359 (.A1(\temp1[4] [20]), .A2(n_1_220), .B1(\temp2[4] [20]), 
      .B2(n_1_219), .C1(n_153), .C2(n_1_218), .ZN(n_1_204));
   INV_X1 i_1_360 (.A(n_1_205), .ZN(n_138));
   AOI222_X1 i_1_361 (.A1(\temp1[4] [21]), .A2(n_1_220), .B1(\temp2[4] [21]), 
      .B2(n_1_219), .C1(n_154), .C2(n_1_218), .ZN(n_1_205));
   INV_X1 i_1_362 (.A(n_1_206), .ZN(n_139));
   AOI222_X1 i_1_363 (.A1(\temp1[4] [22]), .A2(n_1_220), .B1(\temp2[4] [22]), 
      .B2(n_1_219), .C1(n_155), .C2(n_1_218), .ZN(n_1_206));
   INV_X1 i_1_364 (.A(n_1_207), .ZN(n_140));
   AOI222_X1 i_1_365 (.A1(\temp1[4] [23]), .A2(n_1_220), .B1(\temp2[4] [23]), 
      .B2(n_1_219), .C1(n_156), .C2(n_1_218), .ZN(n_1_207));
   INV_X1 i_1_366 (.A(n_1_208), .ZN(n_141));
   AOI222_X1 i_1_367 (.A1(\temp1[4] [24]), .A2(n_1_220), .B1(\temp2[4] [24]), 
      .B2(n_1_219), .C1(n_157), .C2(n_1_218), .ZN(n_1_208));
   INV_X1 i_1_368 (.A(n_1_209), .ZN(n_142));
   AOI222_X1 i_1_369 (.A1(\temp1[4] [25]), .A2(n_1_220), .B1(\temp2[4] [25]), 
      .B2(n_1_219), .C1(n_158), .C2(n_1_218), .ZN(n_1_209));
   INV_X1 i_1_370 (.A(n_1_210), .ZN(n_143));
   AOI222_X1 i_1_371 (.A1(\temp1[4] [26]), .A2(n_1_220), .B1(\temp2[4] [26]), 
      .B2(n_1_219), .C1(n_159), .C2(n_1_218), .ZN(n_1_210));
   INV_X1 i_1_372 (.A(n_1_211), .ZN(n_144));
   AOI222_X1 i_1_373 (.A1(\temp1[4] [27]), .A2(n_1_220), .B1(\temp2[4] [27]), 
      .B2(n_1_219), .C1(n_160), .C2(n_1_218), .ZN(n_1_211));
   INV_X1 i_1_374 (.A(n_1_212), .ZN(n_145));
   AOI222_X1 i_1_375 (.A1(\temp1[4] [28]), .A2(n_1_220), .B1(\temp2[4] [28]), 
      .B2(n_1_219), .C1(n_161), .C2(n_1_218), .ZN(n_1_212));
   INV_X1 i_1_376 (.A(n_1_213), .ZN(n_146));
   AOI222_X1 i_1_377 (.A1(\temp2[4] [29]), .A2(n_1_219), .B1(\temp1[4] [29]), 
      .B2(n_1_220), .C1(n_162), .C2(n_1_218), .ZN(n_1_213));
   INV_X1 i_1_378 (.A(n_1_214), .ZN(n_147));
   AOI222_X1 i_1_379 (.A1(\temp2[4] [30]), .A2(n_1_219), .B1(\temp1[4] [30]), 
      .B2(n_1_220), .C1(n_163), .C2(n_1_218), .ZN(n_1_214));
   INV_X1 i_1_380 (.A(n_1_215), .ZN(n_148));
   AOI221_X1 i_1_381 (.A(n_1_217), .B1(\temp1[4] [31]), .B2(n_1_220), .C1(
      \temp2[4] [31]), .C2(n_1_219), .ZN(n_1_215));
   INV_X1 i_1_382 (.A(n_1_216), .ZN(n_149));
   AOI221_X1 i_1_383 (.A(n_1_217), .B1(\temp1[4] [32]), .B2(n_1_220), .C1(
      \temp2[4] [32]), .C2(n_1_219), .ZN(n_1_216));
   AND2_X1 i_1_384 (.A1(n_164), .A2(n_1_218), .ZN(n_1_217));
   NOR2_X1 i_1_385 (.A1(n_1_220), .A2(n_1_219), .ZN(n_1_218));
   NOR2_X1 i_1_386 (.A1(n_1_18), .A2(r[3]), .ZN(n_1_219));
   NOR2_X1 i_1_387 (.A1(r[4]), .A2(n_1_17), .ZN(n_1_220));
   INV_X1 i_1_388 (.A(n_1_221), .ZN(n_150));
   AOI222_X1 i_1_389 (.A1(\temp1[3] [18]), .A2(n_1_239), .B1(\temp2[3] [18]), 
      .B2(n_1_238), .C1(n_166), .C2(n_1_237), .ZN(n_1_221));
   INV_X1 i_1_390 (.A(n_1_222), .ZN(n_151));
   AOI222_X1 i_1_391 (.A1(\temp2[3] [19]), .A2(n_1_238), .B1(\temp1[3] [19]), 
      .B2(n_1_239), .C1(n_167), .C2(n_1_237), .ZN(n_1_222));
   INV_X1 i_1_392 (.A(n_1_223), .ZN(n_152));
   AOI222_X1 i_1_393 (.A1(\temp2[3] [20]), .A2(n_1_238), .B1(\temp1[3] [20]), 
      .B2(n_1_239), .C1(n_168), .C2(n_1_237), .ZN(n_1_223));
   INV_X1 i_1_394 (.A(n_1_224), .ZN(n_153));
   AOI222_X1 i_1_395 (.A1(\temp2[3] [21]), .A2(n_1_238), .B1(\temp1[3] [21]), 
      .B2(n_1_239), .C1(n_169), .C2(n_1_237), .ZN(n_1_224));
   INV_X1 i_1_396 (.A(n_1_225), .ZN(n_154));
   AOI222_X1 i_1_397 (.A1(\temp2[3] [22]), .A2(n_1_238), .B1(\temp1[3] [22]), 
      .B2(n_1_239), .C1(n_170), .C2(n_1_237), .ZN(n_1_225));
   INV_X1 i_1_398 (.A(n_1_226), .ZN(n_155));
   AOI222_X1 i_1_399 (.A1(\temp2[3] [23]), .A2(n_1_238), .B1(\temp1[3] [23]), 
      .B2(n_1_239), .C1(n_171), .C2(n_1_237), .ZN(n_1_226));
   INV_X1 i_1_400 (.A(n_1_227), .ZN(n_156));
   AOI222_X1 i_1_401 (.A1(\temp2[3] [24]), .A2(n_1_238), .B1(\temp1[3] [24]), 
      .B2(n_1_239), .C1(n_172), .C2(n_1_237), .ZN(n_1_227));
   INV_X1 i_1_402 (.A(n_1_228), .ZN(n_157));
   AOI222_X1 i_1_403 (.A1(\temp2[3] [25]), .A2(n_1_238), .B1(\temp1[3] [25]), 
      .B2(n_1_239), .C1(n_173), .C2(n_1_237), .ZN(n_1_228));
   INV_X1 i_1_404 (.A(n_1_229), .ZN(n_158));
   AOI222_X1 i_1_405 (.A1(\temp2[3] [26]), .A2(n_1_238), .B1(\temp1[3] [26]), 
      .B2(n_1_239), .C1(n_174), .C2(n_1_237), .ZN(n_1_229));
   INV_X1 i_1_406 (.A(n_1_230), .ZN(n_159));
   AOI222_X1 i_1_407 (.A1(\temp2[3] [27]), .A2(n_1_238), .B1(\temp1[3] [27]), 
      .B2(n_1_239), .C1(n_175), .C2(n_1_237), .ZN(n_1_230));
   INV_X1 i_1_408 (.A(n_1_231), .ZN(n_160));
   AOI222_X1 i_1_409 (.A1(\temp2[3] [28]), .A2(n_1_238), .B1(\temp1[3] [28]), 
      .B2(n_1_239), .C1(n_176), .C2(n_1_237), .ZN(n_1_231));
   INV_X1 i_1_410 (.A(n_1_232), .ZN(n_161));
   AOI222_X1 i_1_411 (.A1(\temp2[3] [29]), .A2(n_1_238), .B1(\temp1[3] [29]), 
      .B2(n_1_239), .C1(n_177), .C2(n_1_237), .ZN(n_1_232));
   INV_X1 i_1_412 (.A(n_1_233), .ZN(n_162));
   AOI222_X1 i_1_413 (.A1(\temp2[3] [30]), .A2(n_1_238), .B1(\temp1[3] [30]), 
      .B2(n_1_239), .C1(n_178), .C2(n_1_237), .ZN(n_1_233));
   INV_X1 i_1_414 (.A(n_1_234), .ZN(n_163));
   AOI221_X1 i_1_415 (.A(n_1_236), .B1(\temp1[3] [31]), .B2(n_1_239), .C1(
      \temp2[3] [31]), .C2(n_1_238), .ZN(n_1_234));
   INV_X1 i_1_416 (.A(n_1_235), .ZN(n_164));
   AOI221_X1 i_1_417 (.A(n_1_236), .B1(\temp1[3] [32]), .B2(n_1_239), .C1(
      \temp2[3] [32]), .C2(n_1_238), .ZN(n_1_235));
   AND2_X1 i_1_418 (.A1(n_179), .A2(n_1_237), .ZN(n_1_236));
   NOR2_X1 i_1_419 (.A1(n_1_239), .A2(n_1_238), .ZN(n_1_237));
   NOR2_X1 i_1_420 (.A1(n_1_17), .A2(r[2]), .ZN(n_1_238));
   NOR2_X1 i_1_421 (.A1(r[3]), .A2(n_1_16), .ZN(n_1_239));
   INV_X1 i_1_422 (.A(n_1_240), .ZN(n_165));
   AOI222_X1 i_1_423 (.A1(\temp2[2] [18]), .A2(n_1_257), .B1(\temp1[2] [18]), 
      .B2(n_1_258), .C1(n_181), .C2(n_1_256), .ZN(n_1_240));
   INV_X1 i_1_424 (.A(n_1_241), .ZN(n_166));
   AOI222_X1 i_1_425 (.A1(\temp2[2] [19]), .A2(n_1_257), .B1(\temp1[2] [19]), 
      .B2(n_1_258), .C1(n_182), .C2(n_1_256), .ZN(n_1_241));
   INV_X1 i_1_426 (.A(n_1_242), .ZN(n_167));
   AOI222_X1 i_1_427 (.A1(\temp2[2] [20]), .A2(n_1_257), .B1(\temp1[2] [20]), 
      .B2(n_1_258), .C1(n_183), .C2(n_1_256), .ZN(n_1_242));
   INV_X1 i_1_428 (.A(n_1_243), .ZN(n_168));
   AOI222_X1 i_1_429 (.A1(\temp2[2] [21]), .A2(n_1_257), .B1(\temp1[2] [21]), 
      .B2(n_1_258), .C1(n_184), .C2(n_1_256), .ZN(n_1_243));
   INV_X1 i_1_430 (.A(n_1_244), .ZN(n_169));
   AOI222_X1 i_1_431 (.A1(\temp2[2] [22]), .A2(n_1_257), .B1(\temp1[2] [22]), 
      .B2(n_1_258), .C1(n_185), .C2(n_1_256), .ZN(n_1_244));
   INV_X1 i_1_432 (.A(n_1_245), .ZN(n_170));
   AOI222_X1 i_1_433 (.A1(\temp2[2] [23]), .A2(n_1_257), .B1(\temp1[2] [23]), 
      .B2(n_1_258), .C1(n_186), .C2(n_1_256), .ZN(n_1_245));
   INV_X1 i_1_434 (.A(n_1_246), .ZN(n_171));
   AOI222_X1 i_1_435 (.A1(\temp2[2] [24]), .A2(n_1_257), .B1(\temp1[2] [24]), 
      .B2(n_1_258), .C1(n_187), .C2(n_1_256), .ZN(n_1_246));
   INV_X1 i_1_436 (.A(n_1_247), .ZN(n_172));
   AOI222_X1 i_1_437 (.A1(\temp2[2] [25]), .A2(n_1_257), .B1(\temp1[2] [25]), 
      .B2(n_1_258), .C1(n_188), .C2(n_1_256), .ZN(n_1_247));
   INV_X1 i_1_438 (.A(n_1_248), .ZN(n_173));
   AOI222_X1 i_1_439 (.A1(\temp2[2] [26]), .A2(n_1_257), .B1(\temp1[2] [26]), 
      .B2(n_1_258), .C1(n_189), .C2(n_1_256), .ZN(n_1_248));
   INV_X1 i_1_440 (.A(n_1_249), .ZN(n_174));
   AOI222_X1 i_1_441 (.A1(\temp2[2] [27]), .A2(n_1_257), .B1(\temp1[2] [27]), 
      .B2(n_1_258), .C1(n_190), .C2(n_1_256), .ZN(n_1_249));
   INV_X1 i_1_442 (.A(n_1_250), .ZN(n_175));
   AOI222_X1 i_1_443 (.A1(\temp2[2] [28]), .A2(n_1_257), .B1(\temp1[2] [28]), 
      .B2(n_1_258), .C1(n_191), .C2(n_1_256), .ZN(n_1_250));
   INV_X1 i_1_444 (.A(n_1_251), .ZN(n_176));
   AOI222_X1 i_1_445 (.A1(\temp2[2] [29]), .A2(n_1_257), .B1(\temp1[2] [29]), 
      .B2(n_1_258), .C1(n_192), .C2(n_1_256), .ZN(n_1_251));
   INV_X1 i_1_446 (.A(n_1_252), .ZN(n_177));
   AOI222_X1 i_1_447 (.A1(\temp2[2] [30]), .A2(n_1_257), .B1(\temp1[2] [30]), 
      .B2(n_1_258), .C1(n_193), .C2(n_1_256), .ZN(n_1_252));
   INV_X1 i_1_448 (.A(n_1_253), .ZN(n_178));
   AOI221_X1 i_1_449 (.A(n_1_255), .B1(\temp1[2] [31]), .B2(n_1_258), .C1(
      \temp2[2] [31]), .C2(n_1_257), .ZN(n_1_253));
   INV_X1 i_1_450 (.A(n_1_254), .ZN(n_179));
   AOI221_X1 i_1_451 (.A(n_1_255), .B1(\temp1[2] [32]), .B2(n_1_258), .C1(
      \temp2[2] [32]), .C2(n_1_257), .ZN(n_1_254));
   AND2_X1 i_1_452 (.A1(n_194), .A2(n_1_256), .ZN(n_1_255));
   NOR2_X1 i_1_453 (.A1(n_1_258), .A2(n_1_257), .ZN(n_1_256));
   NOR2_X1 i_1_454 (.A1(n_1_16), .A2(r[1]), .ZN(n_1_257));
   NOR2_X1 i_1_455 (.A1(r[2]), .A2(n_1_15), .ZN(n_1_258));
   INV_X1 i_1_456 (.A(n_1_259), .ZN(n_180));
   AOI222_X1 i_1_457 (.A1(\temp1[1] [18]), .A2(n_1_13), .B1(r[1]), .B2(n_196), 
      .C1(\temp2[1] [18]), .C2(n_1_274), .ZN(n_1_259));
   INV_X1 i_1_458 (.A(n_1_260), .ZN(n_181));
   AOI222_X1 i_1_459 (.A1(mn[3]), .A2(n_1_12), .B1(\temp2[1] [19]), .B2(n_1_274), 
      .C1(\temp1[1] [19]), .C2(n_1_13), .ZN(n_1_260));
   INV_X1 i_1_460 (.A(n_1_261), .ZN(n_182));
   AOI222_X1 i_1_461 (.A1(mn[4]), .A2(n_1_12), .B1(\temp2[1] [20]), .B2(n_1_274), 
      .C1(\temp1[1] [20]), .C2(n_1_13), .ZN(n_1_261));
   INV_X1 i_1_462 (.A(n_1_262), .ZN(n_183));
   AOI222_X1 i_1_463 (.A1(mn[5]), .A2(n_1_12), .B1(\temp2[1] [21]), .B2(n_1_274), 
      .C1(\temp1[1] [21]), .C2(n_1_13), .ZN(n_1_262));
   INV_X1 i_1_464 (.A(n_1_263), .ZN(n_184));
   AOI222_X1 i_1_465 (.A1(mn[6]), .A2(n_1_12), .B1(\temp2[1] [22]), .B2(n_1_274), 
      .C1(\temp1[1] [22]), .C2(n_1_13), .ZN(n_1_263));
   INV_X1 i_1_466 (.A(n_1_264), .ZN(n_185));
   AOI222_X1 i_1_467 (.A1(mn[7]), .A2(n_1_12), .B1(\temp2[1] [23]), .B2(n_1_274), 
      .C1(\temp1[1] [23]), .C2(n_1_13), .ZN(n_1_264));
   INV_X1 i_1_468 (.A(n_1_265), .ZN(n_186));
   AOI222_X1 i_1_469 (.A1(mn[8]), .A2(n_1_12), .B1(\temp2[1] [24]), .B2(n_1_274), 
      .C1(\temp1[1] [24]), .C2(n_1_13), .ZN(n_1_265));
   INV_X1 i_1_470 (.A(n_1_266), .ZN(n_187));
   AOI222_X1 i_1_471 (.A1(mn[9]), .A2(n_1_12), .B1(\temp2[1] [25]), .B2(n_1_274), 
      .C1(\temp1[1] [25]), .C2(n_1_13), .ZN(n_1_266));
   INV_X1 i_1_472 (.A(n_1_267), .ZN(n_188));
   AOI222_X1 i_1_473 (.A1(mn[10]), .A2(n_1_12), .B1(\temp2[1] [26]), .B2(n_1_274), 
      .C1(\temp1[1] [26]), .C2(n_1_13), .ZN(n_1_267));
   INV_X1 i_1_474 (.A(n_1_268), .ZN(n_189));
   AOI222_X1 i_1_475 (.A1(r[1]), .A2(n_205), .B1(\temp2[1] [27]), .B2(n_1_274), 
      .C1(\temp1[1] [27]), .C2(n_1_13), .ZN(n_1_268));
   INV_X1 i_1_476 (.A(n_1_269), .ZN(n_190));
   AOI222_X1 i_1_477 (.A1(r[1]), .A2(n_206), .B1(\temp2[1] [28]), .B2(n_1_274), 
      .C1(\temp1[1] [28]), .C2(n_1_13), .ZN(n_1_269));
   INV_X1 i_1_478 (.A(n_1_270), .ZN(n_191));
   AOI222_X1 i_1_479 (.A1(r[1]), .A2(n_207), .B1(\temp2[1] [29]), .B2(n_1_274), 
      .C1(\temp1[1] [29]), .C2(n_1_13), .ZN(n_1_270));
   INV_X1 i_1_480 (.A(n_1_271), .ZN(n_192));
   AOI222_X1 i_1_481 (.A1(r[1]), .A2(n_208), .B1(\temp2[1] [30]), .B2(n_1_274), 
      .C1(\temp1[1] [30]), .C2(n_1_13), .ZN(n_1_271));
   INV_X1 i_1_482 (.A(n_1_272), .ZN(n_193));
   AOI221_X1 i_1_483 (.A(n_1_275), .B1(\temp2[1] [31]), .B2(n_1_274), .C1(
      \temp1[1] [31]), .C2(n_1_13), .ZN(n_1_272));
   INV_X1 i_1_484 (.A(n_1_273), .ZN(n_194));
   AOI221_X1 i_1_485 (.A(n_1_275), .B1(\temp2[1] [32]), .B2(n_1_274), .C1(
      \temp1[1] [32]), .C2(n_1_13), .ZN(n_1_273));
   NOR2_X1 i_1_486 (.A1(n_1_15), .A2(r[0]), .ZN(n_1_274));
   AND2_X1 i_1_487 (.A1(mn[15]), .A2(n_1_12), .ZN(n_1_275));
   NOR2_X1 i_1_488 (.A1(n_1_15), .A2(n_1_14), .ZN(n_1_12));
   NOR2_X1 i_1_489 (.A1(r[1]), .A2(n_1_14), .ZN(n_1_13));
   AND2_X1 i_1_490 (.A1(r[0]), .A2(mn[1]), .ZN(n_195));
   AND2_X1 i_1_491 (.A1(r[0]), .A2(mn[2]), .ZN(n_196));
   AND2_X1 i_1_492 (.A1(r[0]), .A2(mn[3]), .ZN(n_197));
   AND2_X1 i_1_493 (.A1(r[0]), .A2(mn[4]), .ZN(n_198));
   AND2_X1 i_1_494 (.A1(r[0]), .A2(mn[5]), .ZN(n_199));
   AND2_X1 i_1_495 (.A1(r[0]), .A2(mn[6]), .ZN(n_200));
   AND2_X1 i_1_496 (.A1(r[0]), .A2(mn[7]), .ZN(n_201));
   AND2_X1 i_1_497 (.A1(r[0]), .A2(mn[8]), .ZN(n_202));
   AND2_X1 i_1_498 (.A1(r[0]), .A2(mn[9]), .ZN(n_203));
   AND2_X1 i_1_499 (.A1(r[0]), .A2(mn[10]), .ZN(n_204));
   AND2_X1 i_1_500 (.A1(r[0]), .A2(mn[11]), .ZN(n_205));
   AND2_X1 i_1_501 (.A1(r[0]), .A2(mn[12]), .ZN(n_206));
   AND2_X1 i_1_502 (.A1(r[0]), .A2(mn[13]), .ZN(n_207));
   AND2_X1 i_1_503 (.A1(r[0]), .A2(mn[14]), .ZN(n_208));
   AND2_X1 i_1_504 (.A1(r[0]), .A2(mn[15]), .ZN(n_209));
   INV_X1 i_1_505 (.A(r[0]), .ZN(n_1_14));
   INV_X1 i_1_506 (.A(r[1]), .ZN(n_1_15));
   INV_X1 i_1_507 (.A(r[2]), .ZN(n_1_16));
   INV_X1 i_1_508 (.A(r[3]), .ZN(n_1_17));
   INV_X1 i_1_509 (.A(r[4]), .ZN(n_1_18));
   INV_X1 i_1_510 (.A(r[5]), .ZN(n_1_19));
   INV_X1 i_1_511 (.A(r[6]), .ZN(n_1_20));
   INV_X1 i_1_512 (.A(r[7]), .ZN(n_1_21));
   INV_X1 i_1_513 (.A(r[8]), .ZN(n_1_22));
   INV_X1 i_1_514 (.A(r[9]), .ZN(n_1_23));
   INV_X1 i_1_515 (.A(r[10]), .ZN(n_1_24));
   INV_X1 i_1_516 (.A(r[11]), .ZN(n_1_25));
   INV_X1 i_1_517 (.A(r[12]), .ZN(n_1_26));
   INV_X1 i_1_518 (.A(r[13]), .ZN(n_1_27));
endmodule

module mux__2_5005__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5008__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5011__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5014__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5017__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5020__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5023__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5026__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5029__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5032__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5035__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5038__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5041__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_5044__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__2_0__1(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1__2_2__1(A, B, Cin, sum, overFlow);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output overFlow;

   wire Carry;

   mux__2_5005__1 muxx_1_muxx_j (.sel(B[0]), .in1(), .in2(), .i1(), .i2(B[1]), 
      .out1(sum[1]), .Carry(n_5));
   mux__2_5008__1 muxx_2_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(B[2]), 
      .out1(sum[2]), .Carry(n_9));
   mux__2_5011__1 muxx_3_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(B[3]), 
      .out1(sum[3]), .Carry(n_0));
   mux__2_5014__1 muxx_4_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(B[4]), 
      .out1(sum[4]), .Carry(n_1));
   mux__2_5017__1 muxx_5_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(B[5]), 
      .out1(sum[5]), .Carry(n_2));
   mux__2_5020__1 muxx_6_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(B[6]), 
      .out1(sum[6]), .Carry(n_3));
   mux__2_5023__1 muxx_7_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(B[7]), 
      .out1(sum[7]), .Carry(n_4));
   mux__2_5026__1 muxx_8_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(B[8]), 
      .out1(sum[8]), .Carry(n_6));
   mux__2_5029__1 muxx_9_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(B[9]), 
      .out1(sum[9]), .Carry(n_7));
   mux__2_5032__1 muxx_10_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(B[10]), 
      .out1(sum[10]), .Carry(n_8));
   mux__2_5035__1 muxx_11_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(B[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__2_5038__1 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(B[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__2_5041__1 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(B[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__2_5044__1 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(B[14]), 
      .out1(sum[14]), .Carry(Carry));
   mux__2_0__1 muxx_15_muxx_j (.sel(Carry), .in1(B[15]), .in2(), .i1(), .i2(), 
      .out1(sum[15]), .Carry());
endmodule

module Partial_Full_Adder__2_601__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_597__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_593__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_589__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_585__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_581__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_577__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_573__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_569__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_565__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_561__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_557__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_553__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_549__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_545__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_541__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_634__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_601__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_597__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_593__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_589__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_585__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_581__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_577__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_573__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_569__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_565__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_561__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_557__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_553__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_549__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_545__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_541__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_769__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_765__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_761__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_757__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_753__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_749__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_745__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_741__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_737__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_733__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_729__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_725__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_721__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_717__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_713__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_709__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_802__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_769__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_765__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_761__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_757__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_753__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_749__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_745__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_741__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_737__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_733__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_729__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_725__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_721__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_717__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_713__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_709__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_937__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_933__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_929__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_925__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_921__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_917__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_913__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_909__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_905__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_901__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_897__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_893__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_889__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_885__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_881__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_877__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_970__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_937__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_933__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_929__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_925__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_921__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_917__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_913__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_909__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_905__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_901__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_897__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_893__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_889__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_885__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_881__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_877__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1105__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1101__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1097__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1093__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1089__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1085__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1081__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1077__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1073__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1069__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1065__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1061__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1057__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1053__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1049__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1045__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1138__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1105__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1101__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1097__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1093__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1089__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1085__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1081__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1077__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1073__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1069__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1065__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1061__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1057__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1053__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1049__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1045__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1273__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1269__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1265__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1261__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1257__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1253__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1249__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1245__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1241__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1237__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1233__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1229__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1225__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1221__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1217__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1213__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1306__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1273__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1269__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1265__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1261__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1257__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1253__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1249__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1245__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1241__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1237__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1233__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1229__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1225__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1221__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1217__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1213__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1441__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1437__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1433__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1429__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1425__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1421__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1417__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1413__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1409__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1405__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1401__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1397__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1393__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1389__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1385__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1381__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1474__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1441__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1437__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1433__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1429__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1425__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1421__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1417__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1413__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1409__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1405__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1401__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1397__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1393__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1389__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1385__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1381__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1609__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1605__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1601__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1597__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1593__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1589__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1585__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1581__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1577__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1573__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1569__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1565__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1561__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1557__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1553__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1549__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1642__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1609__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1605__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1601__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1597__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1593__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1589__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1585__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1581__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1577__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1573__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1569__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1565__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1561__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1557__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1553__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1549__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1777__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1773__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1769__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1765__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1761__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1757__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1753__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1749__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1745__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1741__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1737__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1733__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1729__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1725__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1721__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1717__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1810__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1777__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1773__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1769__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1765__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1761__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1757__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1753__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1749__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1745__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1741__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1737__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1733__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1729__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1725__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1721__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1717__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_1945__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_1941__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1937__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1933__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1929__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1925__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1921__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1917__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1913__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1909__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1905__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1901__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1897__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1893__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1889__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_1885__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_1978__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_1945__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_1941__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_1937__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_1933__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_1929__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_1925__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_1921__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_1917__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_1913__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_1909__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_1905__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_1901__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_1897__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_1893__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_1889__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_1885__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2113__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2109__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2105__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2101__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2097__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2093__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2089__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2085__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2081__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2077__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2073__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2069__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2065__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2061__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2057__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2053__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2146__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2113__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2109__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2105__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2101__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2097__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2093__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2089__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2085__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2081__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2077__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2073__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2069__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2065__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2061__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2057__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2053__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2281__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2277__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2273__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2269__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2265__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2261__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2257__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2253__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2249__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2245__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2241__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2237__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2233__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2229__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2225__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2221__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2314__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2281__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2277__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2273__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2269__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2265__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2261__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2257__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2253__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2249__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2245__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2241__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2237__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2233__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2229__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2225__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2221__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2449__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2445__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2441__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2437__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2433__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2429__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2425__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2421__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2417__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2413__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2409__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2405__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2401__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2397__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2393__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2389__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2482__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2449__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2445__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2441__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2437__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2433__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2429__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2425__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2421__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2417__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2413__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2409__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2405__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2401__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2397__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2393__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2389__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2617__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2613__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2609__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2605__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2601__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2597__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2593__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2589__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2585__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2581__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2577__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2573__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2569__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2565__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2561__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2557__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2650__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2617__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2613__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2609__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2605__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2601__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2597__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2593__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2589__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2585__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2581__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2577__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2573__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2569__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2565__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2561__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2557__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2785__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2781__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2777__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2773__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2769__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2765__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2761__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2757__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2753__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2749__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2745__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2741__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2737__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2733__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2729__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2725__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2818__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2785__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2781__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2777__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2773__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2769__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2765__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2761__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2757__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2753__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2749__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2745__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2741__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2737__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2733__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2729__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2725__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_2953__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_2949__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2945__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2941__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2937__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2933__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2929__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2925__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2921__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2917__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2913__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2909__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2905__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2901__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2897__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_2893__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_2986__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_2953__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_2949__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_2945__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_2941__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_2937__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_2933__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_2929__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_2925__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_2921__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_2917__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_2913__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_2909__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_2905__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_2901__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_2897__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_2893__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3121__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3117__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3113__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3109__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3105__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3101__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3097__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3093__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3089__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3085__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3081__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3077__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3073__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3069__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3065__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3061__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3154__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3121__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3117__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3113__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3109__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3105__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3101__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3097__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3093__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3089__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3085__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3081__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3077__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3073__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3069__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3065__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3061__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3289__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3285__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3281__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3277__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3273__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3269__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3265__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3261__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3257__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3253__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3249__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3245__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3241__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3237__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3233__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3229__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3322__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3289__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3285__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3281__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3277__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3273__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3269__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3265__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3261__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3257__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3253__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3249__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3245__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3241__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3237__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3233__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3229__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3457__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3453__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3449__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3445__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3441__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3437__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3433__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3429__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3425__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3421__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3417__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3413__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3409__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3405__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3401__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3397__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3490__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3457__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3453__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3449__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3445__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3441__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3437__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3433__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3429__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3425__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3421__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3417__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3413__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3409__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3405__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3401__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3397__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3625__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3621__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3617__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3613__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3609__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3605__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3601__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3597__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3593__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3589__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3585__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3581__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3577__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3573__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3569__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3565__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3658__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3625__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3621__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3617__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3613__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3609__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3605__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3601__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3597__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3593__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3589__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3585__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3581__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3577__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3573__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3569__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3565__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3793__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3789__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3785__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3781__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3777__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3773__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3769__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3765__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3761__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3757__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3753__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3749__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3745__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3741__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3737__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3733__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3826__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3793__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3789__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3785__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3781__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3777__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3773__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3769__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3765__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3761__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3757__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3753__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3749__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3745__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3741__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3737__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3733__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_3961__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_3957__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3953__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3949__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3945__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3941__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3937__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3933__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3929__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3925__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3921__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3917__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3913__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3909__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3905__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_3901__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_3994__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_3961__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_3957__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_3953__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_3949__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_3945__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_3941__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_3937__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_3933__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_3929__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_3925__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_3921__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_3917__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_3913__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_3909__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_3905__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_3901__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4129__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4125__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4121__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4117__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4113__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4109__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4105__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4101__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4097__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4093__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4089__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4085__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4081__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4077__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4073__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4069__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4162__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4129__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4125__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4121__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4117__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4113__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4109__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4105__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4101__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4097__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4093__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4089__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4085__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4081__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4077__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4073__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4069__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4297__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4293__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4289__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4285__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4281__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4277__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4273__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4269__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4265__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4261__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4257__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4253__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4249__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4245__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4241__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4237__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4330__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4297__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4293__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4289__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4285__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4281__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4277__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4273__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4269__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4265__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4261__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4257__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4253__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4249__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4245__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4241__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4237__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4465__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4461__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4457__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4453__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4449__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4445__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4441__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4437__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4433__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4429__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4425__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4421__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4417__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4413__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4409__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4405__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4498__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4465__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4461__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4457__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4453__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4449__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4445__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4441__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4437__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4433__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4429__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4425__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4421__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4417__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4413__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4409__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4405__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4633__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4629__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4625__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4621__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4617__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4613__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4609__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4605__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4601__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4597__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4593__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4589__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4585__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4581__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4577__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4573__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4666__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4633__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4629__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4625__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4621__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4617__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4613__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4609__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4605__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4601__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4597__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4593__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4589__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4585__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4581__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4577__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4573__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4801__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4797__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4793__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4789__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4785__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4781__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4777__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4773__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4769__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4765__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4761__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4757__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4753__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4749__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4745__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4741__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_4834__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4801__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4797__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4793__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4789__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4785__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4781__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4777__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4773__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4769__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4765__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4761__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4757__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4753__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4749__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4745__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4741__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_4969__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_4965__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4961__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4957__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4953__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4949__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4945__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4941__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4937__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4933__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4929__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4925__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4921__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4917__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4913__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_4909__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__2_5002__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_14;
   wire n_0_1;
   wire n_0_15;
   wire n_0_2;
   wire n_0_16;
   wire n_0_3;
   wire n_0_17;
   wire n_0_4;
   wire n_0_18;
   wire n_0_5;
   wire n_0_19;
   wire n_0_6;
   wire n_0_20;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_4969__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_4965__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_32), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_4961__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_31), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_4957__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_30), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_4953__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_29), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_4949__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_28), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_4945__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_27), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_4941__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(), .S(), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_4937__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(), .S(), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_4933__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(), .S(), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_4929__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(), .S(), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_4925__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(), .S(), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_4921__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(), .S(), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_4917__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(), .S(), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_4913__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(), .S(), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_4909__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_0_14));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_0_14), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_0_15));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_0_15), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_16));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_0_16), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_17));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_0_17), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_0_18));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_0_18), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_0_19));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_0_19), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_0_20));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_0_20), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_27));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_27), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_28));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_28), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_29));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_29), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_30));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_30), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_31));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_31), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_32));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_32), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__2_6__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__2_10__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_14__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_18__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_22__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_26__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_30__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_34__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_38__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_42__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_46__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_50__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_54__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_58__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_62__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__2_66__1(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__1(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_14;
   wire n_0_1;
   wire n_0_15;
   wire n_0_2;
   wire n_0_16;
   wire n_0_3;
   wire n_0_17;
   wire n_0_4;
   wire n_0_18;
   wire n_0_5;
   wire n_0_19;
   wire n_0_6;
   wire n_0_20;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__2_6__1 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__2_10__1 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_32), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__2_14__1 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_31), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__2_18__1 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_30), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__2_22__1 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_29), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__2_26__1 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_28), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__2_30__1 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_27), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__2_34__1 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(), .S(), .P(n_11), .G(n_10));
   Partial_Full_Adder__2_38__1 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(), .S(), .P(n_13), .G(n_12));
   Partial_Full_Adder__2_42__1 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(), .S(), .P(n_15), .G(n_14));
   Partial_Full_Adder__2_46__1 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(), .S(), .P(n_17), .G(n_16));
   Partial_Full_Adder__2_50__1 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(), .S(), .P(n_19), .G(n_18));
   Partial_Full_Adder__2_54__1 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(), .S(), .P(n_21), .G(n_20));
   Partial_Full_Adder__2_58__1 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(), .S(), .P(n_23), .G(n_22));
   Partial_Full_Adder__2_62__1 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(), .S(), .P(n_25), .G(n_24));
   Partial_Full_Adder__2_66__1 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_0_14));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_0_14), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_0_15));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_0_15), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_16));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_0_16), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_17));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_0_17), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_0_18));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_0_18), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_0_19));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_0_19), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_0_20));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_0_20), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_27));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_27), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_28));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_28), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_29));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_29), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_30));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_30), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_31));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_31), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_32));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_32), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module booth_multiplier__1(m, r, result, overflow);
   input [15:0]m;
   input [15:0]r;
   output [15:0]result;
   output overflow;

   wire [15:0]mn;
   wire [32:0]\temp1[1] ;
   wire [32:0]\temp2[1] ;
   wire [32:0]\temp1[2] ;
   wire [32:0]\temp2[2] ;
   wire [32:0]\temp1[3] ;
   wire [32:0]\temp2[3] ;
   wire [32:0]\temp1[4] ;
   wire [32:0]\temp2[4] ;
   wire [32:0]\temp1[5] ;
   wire [32:0]\temp2[5] ;
   wire [32:0]\temp1[6] ;
   wire [32:0]\temp2[6] ;
   wire [32:0]\temp1[7] ;
   wire [32:0]\temp2[7] ;
   wire [32:0]\temp1[8] ;
   wire [32:0]\temp2[8] ;
   wire [32:0]\temp1[9] ;
   wire [32:0]\temp2[9] ;
   wire [32:0]\temp1[10] ;
   wire [32:0]\temp2[10] ;
   wire [32:0]\temp1[11] ;
   wire [32:0]\temp2[11] ;
   wire [32:0]\temp1[12] ;
   wire [32:0]\temp2[12] ;
   wire [32:0]\temp1[13] ;
   wire [32:0]\temp2[13] ;
   wire [32:0]\temp2[14] ;
   wire [32:0]\temp1[14] ;
   wire [15:0]notM;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_177;
   wire n_1_178;
   wire n_1_179;
   wire n_1_180;
   wire n_1_181;
   wire n_1_182;
   wire n_1_183;
   wire n_1_184;
   wire n_1_185;
   wire n_1_186;
   wire n_1_187;
   wire n_1_188;
   wire n_1_189;
   wire n_1_190;
   wire n_1_191;
   wire n_1_192;
   wire n_1_193;
   wire n_1_194;
   wire n_1_195;
   wire n_1_196;
   wire n_1_197;
   wire n_1_198;
   wire n_1_199;
   wire n_1_200;
   wire n_1_201;
   wire n_1_202;
   wire n_1_203;
   wire n_1_204;
   wire n_1_205;
   wire n_1_206;
   wire n_1_207;
   wire n_1_208;
   wire n_1_209;
   wire n_1_210;
   wire n_1_211;
   wire n_1_212;
   wire n_1_213;
   wire n_1_214;
   wire n_1_215;
   wire n_1_216;
   wire n_1_217;
   wire n_1_218;
   wire n_1_219;
   wire n_1_220;
   wire n_1_221;
   wire n_1_222;
   wire n_1_223;
   wire n_1_224;
   wire n_1_225;
   wire n_1_226;
   wire n_1_227;
   wire n_1_228;
   wire n_1_229;
   wire n_1_230;
   wire n_1_231;
   wire n_1_232;
   wire n_1_233;
   wire n_1_234;
   wire n_1_235;
   wire n_1_236;
   wire n_1_237;
   wire n_1_238;
   wire n_1_239;
   wire n_1_240;
   wire n_1_241;
   wire n_1_242;
   wire n_1_243;
   wire n_1_244;
   wire n_1_245;
   wire n_1_246;
   wire n_1_247;
   wire n_1_248;
   wire n_1_249;
   wire n_1_250;
   wire n_1_251;
   wire n_1_252;
   wire n_1_253;
   wire n_1_254;
   wire n_1_255;
   wire n_1_256;
   wire n_1_257;
   wire n_1_258;
   wire n_1_259;
   wire n_1_260;
   wire n_1_261;
   wire n_1_262;
   wire n_1_263;
   wire n_1_264;
   wire n_1_265;
   wire n_1_266;
   wire n_1_267;
   wire n_1_268;
   wire n_1_269;
   wire n_1_270;
   wire n_1_271;
   wire n_1_272;
   wire n_1_273;
   wire n_1_274;
   wire n_1_275;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;

   Addition1__2_2__1 U0 (.A(), .B(notM), .Cin(), .sum({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], uc_0}), .overFlow());
   Carry_Look_Ahead_generic__2_634__1 x_1_Un (.A({n_209, uc_1, n_208, n_207, 
      n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, 
      n_196, n_195, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, 
      uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18}), .B({m[15], m[14], m[13], 
      m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], 
      m[0], uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, 
      uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35}), .Cin(), .S({
      \temp1[1] [32], \temp1[1] [31], \temp1[1] [30], \temp1[1] [29], 
      \temp1[1] [28], \temp1[1] [27], \temp1[1] [26], \temp1[1] [25], 
      \temp1[1] [24], \temp1[1] [23], \temp1[1] [22], \temp1[1] [21], 
      \temp1[1] [20], \temp1[1] [19], \temp1[1] [18], uc_36, uc_37, uc_38, uc_39, 
      uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, 
      uc_50, uc_51, uc_52, uc_53}), .overFlow());
   Carry_Look_Ahead_generic__2_802__1 x_1_Ux (.A({n_209, uc_54, n_208, n_207, 
      n_206, n_205, n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, 
      n_196, n_195, uc_55, uc_56, uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, 
      uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71}), .B({
      mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], 
      mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_72, uc_73, uc_74, uc_75, uc_76, 
      uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, 
      uc_87, uc_88}), .Cin(), .S({\temp2[1] [32], \temp2[1] [31], \temp2[1] [30], 
      \temp2[1] [29], \temp2[1] [28], \temp2[1] [27], \temp2[1] [26], 
      \temp2[1] [25], \temp2[1] [24], \temp2[1] [23], \temp2[1] [22], 
      \temp2[1] [21], \temp2[1] [20], \temp2[1] [19], \temp2[1] [18], uc_89, 
      uc_90, uc_91, uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, uc_98, uc_99, 
      uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, uc_106}), .overFlow());
   Carry_Look_Ahead_generic__2_970__1 x_2_Un (.A({n_194, uc_107, n_193, n_192, 
      n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, 
      n_181, n_180, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, 
      uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, 
      uc_124}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_125, uc_126, uc_127, uc_128, 
      uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, 
      uc_138, uc_139, uc_140, uc_141}), .Cin(), .S({\temp1[2] [32], 
      \temp1[2] [31], \temp1[2] [30], \temp1[2] [29], \temp1[2] [28], 
      \temp1[2] [27], \temp1[2] [26], \temp1[2] [25], \temp1[2] [24], 
      \temp1[2] [23], \temp1[2] [22], \temp1[2] [21], \temp1[2] [20], 
      \temp1[2] [19], \temp1[2] [18], uc_142, uc_143, uc_144, uc_145, uc_146, 
      uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, uc_155, 
      uc_156, uc_157, uc_158, uc_159}), .overFlow());
   Carry_Look_Ahead_generic__2_1138__1 x_2_Ux (.A({n_194, uc_160, n_193, n_192, 
      n_191, n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, 
      n_181, n_180, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, 
      uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, 
      uc_177}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_178, uc_179, 
      uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, uc_186, uc_187, uc_188, 
      uc_189, uc_190, uc_191, uc_192, uc_193, uc_194}), .Cin(), .S({
      \temp2[2] [32], \temp2[2] [31], \temp2[2] [30], \temp2[2] [29], 
      \temp2[2] [28], \temp2[2] [27], \temp2[2] [26], \temp2[2] [25], 
      \temp2[2] [24], \temp2[2] [23], \temp2[2] [22], \temp2[2] [21], 
      \temp2[2] [20], \temp2[2] [19], \temp2[2] [18], uc_195, uc_196, uc_197, 
      uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, uc_204, uc_205, uc_206, 
      uc_207, uc_208, uc_209, uc_210, uc_211, uc_212}), .overFlow());
   Carry_Look_Ahead_generic__2_1306__1 x_3_Un (.A({n_179, uc_213, n_178, n_177, 
      n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
      n_166, n_165, uc_214, uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, 
      uc_221, uc_222, uc_223, uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, 
      uc_230}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_231, uc_232, uc_233, uc_234, 
      uc_235, uc_236, uc_237, uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, 
      uc_244, uc_245, uc_246, uc_247}), .Cin(), .S({\temp1[3] [32], 
      \temp1[3] [31], \temp1[3] [30], \temp1[3] [29], \temp1[3] [28], 
      \temp1[3] [27], \temp1[3] [26], \temp1[3] [25], \temp1[3] [24], 
      \temp1[3] [23], \temp1[3] [22], \temp1[3] [21], \temp1[3] [20], 
      \temp1[3] [19], \temp1[3] [18], uc_248, uc_249, uc_250, uc_251, uc_252, 
      uc_253, uc_254, uc_255, uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, 
      uc_262, uc_263, uc_264, uc_265}), .overFlow());
   Carry_Look_Ahead_generic__2_1474__1 x_3_Ux (.A({n_179, uc_266, n_178, n_177, 
      n_176, n_175, n_174, n_173, n_172, n_171, n_170, n_169, n_168, n_167, 
      n_166, n_165, uc_267, uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, 
      uc_274, uc_275, uc_276, uc_277, uc_278, uc_279, uc_280, uc_281, uc_282, 
      uc_283}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_284, uc_285, 
      uc_286, uc_287, uc_288, uc_289, uc_290, uc_291, uc_292, uc_293, uc_294, 
      uc_295, uc_296, uc_297, uc_298, uc_299, uc_300}), .Cin(), .S({
      \temp2[3] [32], \temp2[3] [31], \temp2[3] [30], \temp2[3] [29], 
      \temp2[3] [28], \temp2[3] [27], \temp2[3] [26], \temp2[3] [25], 
      \temp2[3] [24], \temp2[3] [23], \temp2[3] [22], \temp2[3] [21], 
      \temp2[3] [20], \temp2[3] [19], \temp2[3] [18], uc_301, uc_302, uc_303, 
      uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, 
      uc_313, uc_314, uc_315, uc_316, uc_317, uc_318}), .overFlow());
   Carry_Look_Ahead_generic__2_1642__1 x_4_Un (.A({n_164, uc_319, n_163, n_162, 
      n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, 
      n_151, n_150, uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, 
      uc_327, uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, uc_334, uc_335, 
      uc_336}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_337, uc_338, uc_339, uc_340, 
      uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, uc_348, uc_349, 
      uc_350, uc_351, uc_352, uc_353}), .Cin(), .S({\temp1[4] [32], 
      \temp1[4] [31], \temp1[4] [30], \temp1[4] [29], \temp1[4] [28], 
      \temp1[4] [27], \temp1[4] [26], \temp1[4] [25], \temp1[4] [24], 
      \temp1[4] [23], \temp1[4] [22], \temp1[4] [21], \temp1[4] [20], 
      \temp1[4] [19], \temp1[4] [18], uc_354, uc_355, uc_356, uc_357, uc_358, 
      uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, uc_366, uc_367, 
      uc_368, uc_369, uc_370, uc_371}), .overFlow());
   Carry_Look_Ahead_generic__2_1810__1 x_4_Ux (.A({n_164, uc_372, n_163, n_162, 
      n_161, n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, 
      n_151, n_150, uc_373, uc_374, uc_375, uc_376, uc_377, uc_378, uc_379, 
      uc_380, uc_381, uc_382, uc_383, uc_384, uc_385, uc_386, uc_387, uc_388, 
      uc_389}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_390, uc_391, 
      uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, uc_399, uc_400, 
      uc_401, uc_402, uc_403, uc_404, uc_405, uc_406}), .Cin(), .S({
      \temp2[4] [32], \temp2[4] [31], \temp2[4] [30], \temp2[4] [29], 
      \temp2[4] [28], \temp2[4] [27], \temp2[4] [26], \temp2[4] [25], 
      \temp2[4] [24], \temp2[4] [23], \temp2[4] [22], \temp2[4] [21], 
      \temp2[4] [20], \temp2[4] [19], \temp2[4] [18], uc_407, uc_408, uc_409, 
      uc_410, uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, 
      uc_419, uc_420, uc_421, uc_422, uc_423, uc_424}), .overFlow());
   Carry_Look_Ahead_generic__2_1978__1 x_5_Un (.A({n_149, uc_425, n_148, n_147, 
      n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
      n_136, n_135, uc_426, uc_427, uc_428, uc_429, uc_430, uc_431, uc_432, 
      uc_433, uc_434, uc_435, uc_436, uc_437, uc_438, uc_439, uc_440, uc_441, 
      uc_442}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_443, uc_444, uc_445, uc_446, 
      uc_447, uc_448, uc_449, uc_450, uc_451, uc_452, uc_453, uc_454, uc_455, 
      uc_456, uc_457, uc_458, uc_459}), .Cin(), .S({\temp1[5] [32], 
      \temp1[5] [31], \temp1[5] [30], \temp1[5] [29], \temp1[5] [28], 
      \temp1[5] [27], \temp1[5] [26], \temp1[5] [25], \temp1[5] [24], 
      \temp1[5] [23], \temp1[5] [22], \temp1[5] [21], \temp1[5] [20], 
      \temp1[5] [19], \temp1[5] [18], uc_460, uc_461, uc_462, uc_463, uc_464, 
      uc_465, uc_466, uc_467, uc_468, uc_469, uc_470, uc_471, uc_472, uc_473, 
      uc_474, uc_475, uc_476, uc_477}), .overFlow());
   Carry_Look_Ahead_generic__2_2146__1 x_5_Ux (.A({n_149, uc_478, n_148, n_147, 
      n_146, n_145, n_144, n_143, n_142, n_141, n_140, n_139, n_138, n_137, 
      n_136, n_135, uc_479, uc_480, uc_481, uc_482, uc_483, uc_484, uc_485, 
      uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, uc_492, uc_493, uc_494, 
      uc_495}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_496, uc_497, 
      uc_498, uc_499, uc_500, uc_501, uc_502, uc_503, uc_504, uc_505, uc_506, 
      uc_507, uc_508, uc_509, uc_510, uc_511, uc_512}), .Cin(), .S({
      \temp2[5] [32], \temp2[5] [31], \temp2[5] [30], \temp2[5] [29], 
      \temp2[5] [28], \temp2[5] [27], \temp2[5] [26], \temp2[5] [25], 
      \temp2[5] [24], \temp2[5] [23], \temp2[5] [22], \temp2[5] [21], 
      \temp2[5] [20], \temp2[5] [19], \temp2[5] [18], uc_513, uc_514, uc_515, 
      uc_516, uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, 
      uc_525, uc_526, uc_527, uc_528, uc_529, uc_530}), .overFlow());
   Carry_Look_Ahead_generic__2_2314__1 x_6_Un (.A({n_134, uc_531, n_133, n_132, 
      n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
      n_121, n_120, uc_532, uc_533, uc_534, uc_535, uc_536, uc_537, uc_538, 
      uc_539, uc_540, uc_541, uc_542, uc_543, uc_544, uc_545, uc_546, uc_547, 
      uc_548}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_549, uc_550, uc_551, uc_552, 
      uc_553, uc_554, uc_555, uc_556, uc_557, uc_558, uc_559, uc_560, uc_561, 
      uc_562, uc_563, uc_564, uc_565}), .Cin(), .S({\temp1[6] [32], 
      \temp1[6] [31], \temp1[6] [30], \temp1[6] [29], \temp1[6] [28], 
      \temp1[6] [27], \temp1[6] [26], \temp1[6] [25], \temp1[6] [24], 
      \temp1[6] [23], \temp1[6] [22], \temp1[6] [21], \temp1[6] [20], 
      \temp1[6] [19], \temp1[6] [18], uc_566, uc_567, uc_568, uc_569, uc_570, 
      uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, 
      uc_580, uc_581, uc_582, uc_583}), .overFlow());
   Carry_Look_Ahead_generic__2_2482__1 x_6_Ux (.A({n_134, uc_584, n_133, n_132, 
      n_131, n_130, n_129, n_128, n_127, n_126, n_125, n_124, n_123, n_122, 
      n_121, n_120, uc_585, uc_586, uc_587, uc_588, uc_589, uc_590, uc_591, 
      uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, uc_599, uc_600, 
      uc_601}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_602, uc_603, 
      uc_604, uc_605, uc_606, uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, 
      uc_613, uc_614, uc_615, uc_616, uc_617, uc_618}), .Cin(), .S({
      \temp2[6] [32], \temp2[6] [31], \temp2[6] [30], \temp2[6] [29], 
      \temp2[6] [28], \temp2[6] [27], \temp2[6] [26], \temp2[6] [25], 
      \temp2[6] [24], \temp2[6] [23], \temp2[6] [22], \temp2[6] [21], 
      \temp2[6] [20], \temp2[6] [19], \temp2[6] [18], uc_619, uc_620, uc_621, 
      uc_622, uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, uc_629, uc_630, 
      uc_631, uc_632, uc_633, uc_634, uc_635, uc_636}), .overFlow());
   Carry_Look_Ahead_generic__2_2650__1 x_7_Un (.A({n_119, uc_637, n_118, n_117, 
      n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
      n_106, n_105, uc_638, uc_639, uc_640, uc_641, uc_642, uc_643, uc_644, 
      uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, uc_651, uc_652, uc_653, 
      uc_654}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_655, uc_656, uc_657, uc_658, 
      uc_659, uc_660, uc_661, uc_662, uc_663, uc_664, uc_665, uc_666, uc_667, 
      uc_668, uc_669, uc_670, uc_671}), .Cin(), .S({\temp1[7] [32], 
      \temp1[7] [31], \temp1[7] [30], \temp1[7] [29], \temp1[7] [28], 
      \temp1[7] [27], \temp1[7] [26], \temp1[7] [25], \temp1[7] [24], 
      \temp1[7] [23], \temp1[7] [22], \temp1[7] [21], \temp1[7] [20], 
      \temp1[7] [19], \temp1[7] [18], uc_672, uc_673, uc_674, uc_675, uc_676, 
      uc_677, uc_678, uc_679, uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, 
      uc_686, uc_687, uc_688, uc_689}), .overFlow());
   Carry_Look_Ahead_generic__2_2818__1 x_7_Ux (.A({n_119, uc_690, n_118, n_117, 
      n_116, n_115, n_114, n_113, n_112, n_111, n_110, n_109, n_108, n_107, 
      n_106, n_105, uc_691, uc_692, uc_693, uc_694, uc_695, uc_696, uc_697, 
      uc_698, uc_699, uc_700, uc_701, uc_702, uc_703, uc_704, uc_705, uc_706, 
      uc_707}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], 
      mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_708, uc_709, 
      uc_710, uc_711, uc_712, uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, 
      uc_719, uc_720, uc_721, uc_722, uc_723, uc_724}), .Cin(), .S({
      \temp2[7] [32], \temp2[7] [31], \temp2[7] [30], \temp2[7] [29], 
      \temp2[7] [28], \temp2[7] [27], \temp2[7] [26], \temp2[7] [25], 
      \temp2[7] [24], \temp2[7] [23], \temp2[7] [22], \temp2[7] [21], 
      \temp2[7] [20], \temp2[7] [19], \temp2[7] [18], uc_725, uc_726, uc_727, 
      uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, uc_734, uc_735, uc_736, 
      uc_737, uc_738, uc_739, uc_740, uc_741, uc_742}), .overFlow());
   Carry_Look_Ahead_generic__2_2986__1 x_8_Un (.A({n_104, uc_743, n_103, n_102, 
      n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
      uc_744, uc_745, uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, 
      uc_753, uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, uc_760}), .B({
      m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_761, uc_762, uc_763, uc_764, uc_765, 
      uc_766, uc_767, uc_768, uc_769, uc_770, uc_771, uc_772, uc_773, uc_774, 
      uc_775, uc_776, uc_777}), .Cin(), .S({\temp1[8] [32], \temp1[8] [31], 
      \temp1[8] [30], \temp1[8] [29], \temp1[8] [28], \temp1[8] [27], 
      \temp1[8] [26], \temp1[8] [25], \temp1[8] [24], \temp1[8] [23], 
      \temp1[8] [22], \temp1[8] [21], \temp1[8] [20], \temp1[8] [19], 
      \temp1[8] [18], uc_778, uc_779, uc_780, uc_781, uc_782, uc_783, uc_784, 
      uc_785, uc_786, uc_787, uc_788, uc_789, uc_790, uc_791, uc_792, uc_793, 
      uc_794, uc_795}), .overFlow());
   Carry_Look_Ahead_generic__2_3154__1 x_8_Ux (.A({n_104, uc_796, n_103, n_102, 
      n_101, n_100, n_99, n_98, n_97, n_96, n_95, n_94, n_93, n_92, n_91, n_90, 
      uc_797, uc_798, uc_799, uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, 
      uc_806, uc_807, uc_808, uc_809, uc_810, uc_811, uc_812, uc_813}), .B({
      mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], 
      mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_814, uc_815, uc_816, uc_817, 
      uc_818, uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, uc_826, 
      uc_827, uc_828, uc_829, uc_830}), .Cin(), .S({\temp2[8] [32], 
      \temp2[8] [31], \temp2[8] [30], \temp2[8] [29], \temp2[8] [28], 
      \temp2[8] [27], \temp2[8] [26], \temp2[8] [25], \temp2[8] [24], 
      \temp2[8] [23], \temp2[8] [22], \temp2[8] [21], \temp2[8] [20], 
      \temp2[8] [19], \temp2[8] [18], uc_831, uc_832, uc_833, uc_834, uc_835, 
      uc_836, uc_837, uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, uc_844, 
      uc_845, uc_846, uc_847, uc_848}), .overFlow());
   Carry_Look_Ahead_generic__2_3322__1 x_9_Un (.A({n_89, uc_849, n_88, n_87, 
      n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, 
      uc_850, uc_851, uc_852, uc_853, uc_854, uc_855, uc_856, uc_857, uc_858, 
      uc_859, uc_860, uc_861, uc_862, uc_863, uc_864, uc_865, uc_866}), .B({
      m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_867, uc_868, uc_869, uc_870, uc_871, 
      uc_872, uc_873, uc_874, uc_875, uc_876, uc_877, uc_878, uc_879, uc_880, 
      uc_881, uc_882, uc_883}), .Cin(), .S({\temp1[9] [32], \temp1[9] [31], 
      \temp1[9] [30], \temp1[9] [29], \temp1[9] [28], \temp1[9] [27], 
      \temp1[9] [26], \temp1[9] [25], \temp1[9] [24], \temp1[9] [23], 
      \temp1[9] [22], \temp1[9] [21], \temp1[9] [20], \temp1[9] [19], 
      \temp1[9] [18], uc_884, uc_885, uc_886, uc_887, uc_888, uc_889, uc_890, 
      uc_891, uc_892, uc_893, uc_894, uc_895, uc_896, uc_897, uc_898, uc_899, 
      uc_900, uc_901}), .overFlow());
   Carry_Look_Ahead_generic__2_3490__1 x_9_Ux (.A({n_89, uc_902, n_88, n_87, 
      n_86, n_85, n_84, n_83, n_82, n_81, n_80, n_79, n_78, n_77, n_76, n_75, 
      uc_903, uc_904, uc_905, uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, 
      uc_912, uc_913, uc_914, uc_915, uc_916, uc_917, uc_918, uc_919}), .B({
      mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], 
      mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_920, uc_921, uc_922, uc_923, 
      uc_924, uc_925, uc_926, uc_927, uc_928, uc_929, uc_930, uc_931, uc_932, 
      uc_933, uc_934, uc_935, uc_936}), .Cin(), .S({\temp2[9] [32], 
      \temp2[9] [31], \temp2[9] [30], \temp2[9] [29], \temp2[9] [28], 
      \temp2[9] [27], \temp2[9] [26], \temp2[9] [25], \temp2[9] [24], 
      \temp2[9] [23], \temp2[9] [22], \temp2[9] [21], \temp2[9] [20], 
      \temp2[9] [19], \temp2[9] [18], uc_937, uc_938, uc_939, uc_940, uc_941, 
      uc_942, uc_943, uc_944, uc_945, uc_946, uc_947, uc_948, uc_949, uc_950, 
      uc_951, uc_952, uc_953, uc_954}), .overFlow());
   Carry_Look_Ahead_generic__2_3658__1 x_10_Un (.A({n_74, uc_955, n_73, n_72, 
      n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
      uc_956, uc_957, uc_958, uc_959, uc_960, uc_961, uc_962, uc_963, uc_964, 
      uc_965, uc_966, uc_967, uc_968, uc_969, uc_970, uc_971, uc_972}), .B({
      m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_973, uc_974, uc_975, uc_976, uc_977, 
      uc_978, uc_979, uc_980, uc_981, uc_982, uc_983, uc_984, uc_985, uc_986, 
      uc_987, uc_988, uc_989}), .Cin(), .S({\temp1[10] [32], \temp1[10] [31], 
      \temp1[10] [30], \temp1[10] [29], \temp1[10] [28], \temp1[10] [27], 
      \temp1[10] [26], \temp1[10] [25], \temp1[10] [24], \temp1[10] [23], 
      \temp1[10] [22], \temp1[10] [21], \temp1[10] [20], \temp1[10] [19], 
      \temp1[10] [18], uc_990, uc_991, uc_992, uc_993, uc_994, uc_995, uc_996, 
      uc_997, uc_998, uc_999, uc_1000, uc_1001, uc_1002, uc_1003, uc_1004, 
      uc_1005, uc_1006, uc_1007}), .overFlow());
   Carry_Look_Ahead_generic__2_3826__1 x_10_Ux (.A({n_74, uc_1008, n_73, n_72, 
      n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64, n_63, n_62, n_61, n_60, 
      uc_1009, uc_1010, uc_1011, uc_1012, uc_1013, uc_1014, uc_1015, uc_1016, 
      uc_1017, uc_1018, uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, uc_1024, 
      uc_1025}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], 
      mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1026, 
      uc_1027, uc_1028, uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, uc_1034, 
      uc_1035, uc_1036, uc_1037, uc_1038, uc_1039, uc_1040, uc_1041, uc_1042}), 
      .Cin(), .S({\temp2[10] [32], \temp2[10] [31], \temp2[10] [30], 
      \temp2[10] [29], \temp2[10] [28], \temp2[10] [27], \temp2[10] [26], 
      \temp2[10] [25], \temp2[10] [24], \temp2[10] [23], \temp2[10] [22], 
      \temp2[10] [21], \temp2[10] [20], \temp2[10] [19], \temp2[10] [18], 
      uc_1043, uc_1044, uc_1045, uc_1046, uc_1047, uc_1048, uc_1049, uc_1050, 
      uc_1051, uc_1052, uc_1053, uc_1054, uc_1055, uc_1056, uc_1057, uc_1058, 
      uc_1059, uc_1060}), .overFlow());
   Carry_Look_Ahead_generic__2_3994__1 x_11_Un (.A({n_59, uc_1061, n_58, n_57, 
      n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, 
      uc_1062, uc_1063, uc_1064, uc_1065, uc_1066, uc_1067, uc_1068, uc_1069, 
      uc_1070, uc_1071, uc_1072, uc_1073, uc_1074, uc_1075, uc_1076, uc_1077, 
      uc_1078}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_1079, uc_1080, uc_1081, 
      uc_1082, uc_1083, uc_1084, uc_1085, uc_1086, uc_1087, uc_1088, uc_1089, 
      uc_1090, uc_1091, uc_1092, uc_1093, uc_1094, uc_1095}), .Cin(), .S({
      \temp1[11] [32], \temp1[11] [31], \temp1[11] [30], \temp1[11] [29], 
      \temp1[11] [28], \temp1[11] [27], \temp1[11] [26], \temp1[11] [25], 
      \temp1[11] [24], \temp1[11] [23], \temp1[11] [22], \temp1[11] [21], 
      \temp1[11] [20], \temp1[11] [19], \temp1[11] [18], uc_1096, uc_1097, 
      uc_1098, uc_1099, uc_1100, uc_1101, uc_1102, uc_1103, uc_1104, uc_1105, 
      uc_1106, uc_1107, uc_1108, uc_1109, uc_1110, uc_1111, uc_1112, uc_1113}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_4162__1 x_11_Ux (.A({n_59, uc_1114, n_58, n_57, 
      n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, 
      uc_1115, uc_1116, uc_1117, uc_1118, uc_1119, uc_1120, uc_1121, uc_1122, 
      uc_1123, uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, uc_1130, 
      uc_1131}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], 
      mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1132, 
      uc_1133, uc_1134, uc_1135, uc_1136, uc_1137, uc_1138, uc_1139, uc_1140, 
      uc_1141, uc_1142, uc_1143, uc_1144, uc_1145, uc_1146, uc_1147, uc_1148}), 
      .Cin(), .S({\temp2[11] [32], \temp2[11] [31], \temp2[11] [30], 
      \temp2[11] [29], \temp2[11] [28], \temp2[11] [27], \temp2[11] [26], 
      \temp2[11] [25], \temp2[11] [24], \temp2[11] [23], \temp2[11] [22], 
      \temp2[11] [21], \temp2[11] [20], \temp2[11] [19], \temp2[11] [18], 
      uc_1149, uc_1150, uc_1151, uc_1152, uc_1153, uc_1154, uc_1155, uc_1156, 
      uc_1157, uc_1158, uc_1159, uc_1160, uc_1161, uc_1162, uc_1163, uc_1164, 
      uc_1165, uc_1166}), .overFlow());
   Carry_Look_Ahead_generic__2_4330__1 x_12_Un (.A({n_44, uc_1167, n_43, n_42, 
      n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
      uc_1168, uc_1169, uc_1170, uc_1171, uc_1172, uc_1173, uc_1174, uc_1175, 
      uc_1176, uc_1177, uc_1178, uc_1179, uc_1180, uc_1181, uc_1182, uc_1183, 
      uc_1184}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_1185, uc_1186, uc_1187, 
      uc_1188, uc_1189, uc_1190, uc_1191, uc_1192, uc_1193, uc_1194, uc_1195, 
      uc_1196, uc_1197, uc_1198, uc_1199, uc_1200, uc_1201}), .Cin(), .S({
      \temp1[12] [32], \temp1[12] [31], \temp1[12] [30], \temp1[12] [29], 
      \temp1[12] [28], \temp1[12] [27], \temp1[12] [26], \temp1[12] [25], 
      \temp1[12] [24], \temp1[12] [23], \temp1[12] [22], \temp1[12] [21], 
      \temp1[12] [20], \temp1[12] [19], \temp1[12] [18], uc_1202, uc_1203, 
      uc_1204, uc_1205, uc_1206, uc_1207, uc_1208, uc_1209, uc_1210, uc_1211, 
      uc_1212, uc_1213, uc_1214, uc_1215, uc_1216, uc_1217, uc_1218, uc_1219}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_4498__1 x_12_Ux (.A({n_44, uc_1220, n_43, n_42, 
      n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, 
      uc_1221, uc_1222, uc_1223, uc_1224, uc_1225, uc_1226, uc_1227, uc_1228, 
      uc_1229, uc_1230, uc_1231, uc_1232, uc_1233, uc_1234, uc_1235, uc_1236, 
      uc_1237}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], 
      mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1238, 
      uc_1239, uc_1240, uc_1241, uc_1242, uc_1243, uc_1244, uc_1245, uc_1246, 
      uc_1247, uc_1248, uc_1249, uc_1250, uc_1251, uc_1252, uc_1253, uc_1254}), 
      .Cin(), .S({\temp2[12] [32], \temp2[12] [31], \temp2[12] [30], 
      \temp2[12] [29], \temp2[12] [28], \temp2[12] [27], \temp2[12] [26], 
      \temp2[12] [25], \temp2[12] [24], \temp2[12] [23], \temp2[12] [22], 
      \temp2[12] [21], \temp2[12] [20], \temp2[12] [19], \temp2[12] [18], 
      uc_1255, uc_1256, uc_1257, uc_1258, uc_1259, uc_1260, uc_1261, uc_1262, 
      uc_1263, uc_1264, uc_1265, uc_1266, uc_1267, uc_1268, uc_1269, uc_1270, 
      uc_1271, uc_1272}), .overFlow());
   Carry_Look_Ahead_generic__2_4666__1 x_13_Un (.A({n_29, uc_1273, n_28, n_27, 
      n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, 
      uc_1274, uc_1275, uc_1276, uc_1277, uc_1278, uc_1279, uc_1280, uc_1281, 
      uc_1282, uc_1283, uc_1284, uc_1285, uc_1286, uc_1287, uc_1288, uc_1289, 
      uc_1290}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], 
      m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_1291, uc_1292, uc_1293, 
      uc_1294, uc_1295, uc_1296, uc_1297, uc_1298, uc_1299, uc_1300, uc_1301, 
      uc_1302, uc_1303, uc_1304, uc_1305, uc_1306, uc_1307}), .Cin(), .S({
      \temp1[13] [32], \temp1[13] [31], \temp1[13] [30], \temp1[13] [29], 
      \temp1[13] [28], \temp1[13] [27], \temp1[13] [26], \temp1[13] [25], 
      \temp1[13] [24], \temp1[13] [23], \temp1[13] [22], \temp1[13] [21], 
      \temp1[13] [20], \temp1[13] [19], \temp1[13] [18], uc_1308, uc_1309, 
      uc_1310, uc_1311, uc_1312, uc_1313, uc_1314, uc_1315, uc_1316, uc_1317, 
      uc_1318, uc_1319, uc_1320, uc_1321, uc_1322, uc_1323, uc_1324, uc_1325}), 
      .overFlow());
   Carry_Look_Ahead_generic__2_4834__1 x_13_Ux (.A({n_29, uc_1326, n_28, n_27, 
      n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16, n_15, 
      uc_1327, uc_1328, uc_1329, uc_1330, uc_1331, uc_1332, uc_1333, uc_1334, 
      uc_1335, uc_1336, uc_1337, uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, 
      uc_1343}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], 
      mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1344, 
      uc_1345, uc_1346, uc_1347, uc_1348, uc_1349, uc_1350, uc_1351, uc_1352, 
      uc_1353, uc_1354, uc_1355, uc_1356, uc_1357, uc_1358, uc_1359, uc_1360}), 
      .Cin(), .S({\temp2[13] [32], \temp2[13] [31], \temp2[13] [30], 
      \temp2[13] [29], \temp2[13] [28], \temp2[13] [27], \temp2[13] [26], 
      \temp2[13] [25], \temp2[13] [24], \temp2[13] [23], \temp2[13] [22], 
      \temp2[13] [21], \temp2[13] [20], \temp2[13] [19], \temp2[13] [18], 
      uc_1361, uc_1362, uc_1363, uc_1364, uc_1365, uc_1366, uc_1367, uc_1368, 
      uc_1369, uc_1370, uc_1371, uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, 
      uc_1377, uc_1378}), .overFlow());
   Carry_Look_Ahead_generic__2_5002__1 x_14_Ux (.A({n_14, uc_1379, n_13, n_12, 
      n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_1380, 
      uc_1381, uc_1382, uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, uc_1388, 
      uc_1389, uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396}), 
      .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], 
      mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_1397, uc_1398, uc_1399, 
      uc_1400, uc_1401, uc_1402, uc_1403, uc_1404, uc_1405, uc_1406, uc_1407, 
      uc_1408, uc_1409, uc_1410, uc_1411, uc_1412, uc_1413}), .Cin(), .S({
      \temp2[14] [32], \temp2[14] [31], \temp2[14] [30], \temp2[14] [29], 
      \temp2[14] [28], \temp2[14] [27], \temp2[14] [26], uc_1414, uc_1415, 
      uc_1416, uc_1417, uc_1418, uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, 
      uc_1424, uc_1425, uc_1426, uc_1427, uc_1428, uc_1429, uc_1430, uc_1431, 
      uc_1432, uc_1433, uc_1434, uc_1435, uc_1436, uc_1437, uc_1438, uc_1439}), 
      .overFlow());
   Carry_Look_Ahead_generic__1 x_14_Un (.A({n_14, uc_1440, n_13, n_12, n_11, 
      n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0, uc_1441, uc_1442, 
      uc_1443, uc_1444, uc_1445, uc_1446, uc_1447, uc_1448, uc_1449, uc_1450, 
      uc_1451, uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, uc_1457}), .B({m[15], 
      m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], 
      m[3], m[2], m[1], m[0], uc_1458, uc_1459, uc_1460, uc_1461, uc_1462, 
      uc_1463, uc_1464, uc_1465, uc_1466, uc_1467, uc_1468, uc_1469, uc_1470, 
      uc_1471, uc_1472, uc_1473, uc_1474}), .Cin(), .S({\temp1[14] [32], 
      \temp1[14] [31], \temp1[14] [30], \temp1[14] [29], \temp1[14] [28], 
      \temp1[14] [27], \temp1[14] [26], uc_1475, uc_1476, uc_1477, uc_1478, 
      uc_1479, uc_1480, uc_1481, uc_1482, uc_1483, uc_1484, uc_1485, uc_1486, 
      uc_1487, uc_1488, uc_1489, uc_1490, uc_1491, uc_1492, uc_1493, uc_1494, 
      uc_1495, uc_1496, uc_1497, uc_1498, uc_1499, uc_1500}), .overFlow());
   INV_X1 i_0_0 (.A(m[0]), .ZN(notM[0]));
   INV_X1 i_0_1 (.A(m[1]), .ZN(notM[1]));
   INV_X1 i_0_2 (.A(m[2]), .ZN(notM[2]));
   INV_X1 i_0_3 (.A(m[3]), .ZN(notM[3]));
   INV_X1 i_0_4 (.A(m[4]), .ZN(notM[4]));
   INV_X1 i_0_5 (.A(m[5]), .ZN(notM[5]));
   INV_X1 i_0_6 (.A(m[6]), .ZN(notM[6]));
   INV_X1 i_0_7 (.A(m[7]), .ZN(notM[7]));
   INV_X1 i_0_8 (.A(m[8]), .ZN(notM[8]));
   INV_X1 i_0_9 (.A(m[9]), .ZN(notM[9]));
   INV_X1 i_0_10 (.A(m[10]), .ZN(notM[10]));
   INV_X1 i_0_11 (.A(m[11]), .ZN(notM[11]));
   INV_X1 i_0_12 (.A(m[12]), .ZN(notM[12]));
   INV_X1 i_0_13 (.A(m[13]), .ZN(notM[13]));
   INV_X1 i_0_14 (.A(m[14]), .ZN(notM[14]));
   INV_X1 i_0_15 (.A(m[15]), .ZN(notM[15]));
   AOI22_X1 i_1_0 (.A1(n_1_3), .A2(n_1_2), .B1(n_1_1), .B2(n_1_0), .ZN(overflow));
   NOR3_X1 i_1_1 (.A1(n_1_9), .A2(n_1_4), .A3(n_1_5), .ZN(n_1_0));
   NOR4_X1 i_1_2 (.A1(n_1_11), .A2(n_1_6), .A3(n_1_8), .A4(n_1_7), .ZN(n_1_1));
   AND3_X1 i_1_3 (.A1(n_1_9), .A2(n_1_7), .A3(n_1_6), .ZN(n_1_2));
   AND4_X1 i_1_4 (.A1(n_1_8), .A2(n_1_4), .A3(n_1_11), .A4(n_1_5), .ZN(n_1_3));
   AOI222_X1 i_1_5 (.A1(\temp1[14] [28]), .A2(n_1_30), .B1(\temp2[14] [28]), 
      .B2(n_1_29), .C1(n_11), .C2(n_1_28), .ZN(n_1_4));
   AOI222_X1 i_1_6 (.A1(\temp1[14] [27]), .A2(n_1_30), .B1(\temp2[14] [27]), 
      .B2(n_1_29), .C1(n_10), .C2(n_1_28), .ZN(n_1_5));
   AOI222_X1 i_1_7 (.A1(\temp1[14] [30]), .A2(n_1_30), .B1(\temp2[14] [30]), 
      .B2(n_1_29), .C1(n_13), .C2(n_1_28), .ZN(n_1_6));
   AOI222_X1 i_1_8 (.A1(\temp1[14] [29]), .A2(n_1_30), .B1(\temp2[14] [29]), 
      .B2(n_1_29), .C1(n_12), .C2(n_1_28), .ZN(n_1_7));
   AOI221_X1 i_1_9 (.A(n_1_10), .B1(\temp1[14] [31]), .B2(n_1_30), .C1(
      \temp2[14] [31]), .C2(n_1_29), .ZN(n_1_8));
   AOI221_X1 i_1_10 (.A(n_1_10), .B1(\temp1[14] [32]), .B2(n_1_30), .C1(
      \temp2[14] [32]), .C2(n_1_29), .ZN(n_1_9));
   AND2_X1 i_1_11 (.A1(n_14), .A2(n_1_28), .ZN(n_1_10));
   AOI222_X1 i_1_12 (.A1(\temp1[14] [26]), .A2(n_1_30), .B1(\temp2[14] [26]), 
      .B2(n_1_29), .C1(n_9), .C2(n_1_28), .ZN(n_1_11));
   NOR2_X1 i_1_45 (.A1(n_1_30), .A2(n_1_29), .ZN(n_1_28));
   AND2_X1 i_1_46 (.A1(r[14]), .A2(n_1_27), .ZN(n_1_29));
   NOR2_X1 i_1_47 (.A1(r[14]), .A2(n_1_27), .ZN(n_1_30));
   INV_X1 i_1_48 (.A(n_1_31), .ZN(n_0));
   AOI222_X1 i_1_49 (.A1(\temp1[13] [18]), .A2(n_1_49), .B1(\temp2[13] [18]), 
      .B2(n_1_48), .C1(n_16), .C2(n_1_47), .ZN(n_1_31));
   INV_X1 i_1_50 (.A(n_1_32), .ZN(n_1));
   AOI222_X1 i_1_51 (.A1(\temp1[13] [19]), .A2(n_1_49), .B1(\temp2[13] [19]), 
      .B2(n_1_48), .C1(n_17), .C2(n_1_47), .ZN(n_1_32));
   INV_X1 i_1_52 (.A(n_1_33), .ZN(n_2));
   AOI222_X1 i_1_53 (.A1(\temp1[13] [20]), .A2(n_1_49), .B1(\temp2[13] [20]), 
      .B2(n_1_48), .C1(n_18), .C2(n_1_47), .ZN(n_1_33));
   INV_X1 i_1_54 (.A(n_1_34), .ZN(n_3));
   AOI222_X1 i_1_55 (.A1(\temp1[13] [21]), .A2(n_1_49), .B1(\temp2[13] [21]), 
      .B2(n_1_48), .C1(n_19), .C2(n_1_47), .ZN(n_1_34));
   INV_X1 i_1_56 (.A(n_1_35), .ZN(n_4));
   AOI222_X1 i_1_57 (.A1(\temp1[13] [22]), .A2(n_1_49), .B1(\temp2[13] [22]), 
      .B2(n_1_48), .C1(n_20), .C2(n_1_47), .ZN(n_1_35));
   INV_X1 i_1_58 (.A(n_1_36), .ZN(n_5));
   AOI222_X1 i_1_59 (.A1(\temp1[13] [23]), .A2(n_1_49), .B1(\temp2[13] [23]), 
      .B2(n_1_48), .C1(n_21), .C2(n_1_47), .ZN(n_1_36));
   INV_X1 i_1_60 (.A(n_1_37), .ZN(n_6));
   AOI222_X1 i_1_61 (.A1(\temp1[13] [24]), .A2(n_1_49), .B1(\temp2[13] [24]), 
      .B2(n_1_48), .C1(n_22), .C2(n_1_47), .ZN(n_1_37));
   INV_X1 i_1_62 (.A(n_1_38), .ZN(n_7));
   AOI222_X1 i_1_63 (.A1(\temp1[13] [25]), .A2(n_1_49), .B1(\temp2[13] [25]), 
      .B2(n_1_48), .C1(n_23), .C2(n_1_47), .ZN(n_1_38));
   INV_X1 i_1_64 (.A(n_1_39), .ZN(n_8));
   AOI222_X1 i_1_65 (.A1(\temp1[13] [26]), .A2(n_1_49), .B1(\temp2[13] [26]), 
      .B2(n_1_48), .C1(n_24), .C2(n_1_47), .ZN(n_1_39));
   INV_X1 i_1_66 (.A(n_1_40), .ZN(n_9));
   AOI222_X1 i_1_67 (.A1(\temp1[13] [27]), .A2(n_1_49), .B1(\temp2[13] [27]), 
      .B2(n_1_48), .C1(n_25), .C2(n_1_47), .ZN(n_1_40));
   INV_X1 i_1_68 (.A(n_1_41), .ZN(n_10));
   AOI222_X1 i_1_69 (.A1(\temp1[13] [28]), .A2(n_1_49), .B1(\temp2[13] [28]), 
      .B2(n_1_48), .C1(n_26), .C2(n_1_47), .ZN(n_1_41));
   INV_X1 i_1_70 (.A(n_1_42), .ZN(n_11));
   AOI222_X1 i_1_71 (.A1(\temp1[13] [29]), .A2(n_1_49), .B1(\temp2[13] [29]), 
      .B2(n_1_48), .C1(n_27), .C2(n_1_47), .ZN(n_1_42));
   INV_X1 i_1_72 (.A(n_1_43), .ZN(n_12));
   AOI222_X1 i_1_73 (.A1(\temp1[13] [30]), .A2(n_1_49), .B1(\temp2[13] [30]), 
      .B2(n_1_48), .C1(n_28), .C2(n_1_47), .ZN(n_1_43));
   INV_X1 i_1_74 (.A(n_1_44), .ZN(n_13));
   AOI221_X1 i_1_75 (.A(n_1_46), .B1(\temp1[13] [31]), .B2(n_1_49), .C1(
      \temp2[13] [31]), .C2(n_1_48), .ZN(n_1_44));
   INV_X1 i_1_76 (.A(n_1_45), .ZN(n_14));
   AOI221_X1 i_1_77 (.A(n_1_46), .B1(\temp1[13] [32]), .B2(n_1_49), .C1(
      \temp2[13] [32]), .C2(n_1_48), .ZN(n_1_45));
   AND2_X1 i_1_78 (.A1(n_29), .A2(n_1_47), .ZN(n_1_46));
   NOR2_X1 i_1_79 (.A1(n_1_49), .A2(n_1_48), .ZN(n_1_47));
   NOR2_X1 i_1_80 (.A1(n_1_27), .A2(r[12]), .ZN(n_1_48));
   NOR2_X1 i_1_81 (.A1(r[13]), .A2(n_1_26), .ZN(n_1_49));
   INV_X1 i_1_82 (.A(n_1_50), .ZN(n_15));
   AOI222_X1 i_1_83 (.A1(\temp1[12] [18]), .A2(n_1_68), .B1(\temp2[12] [18]), 
      .B2(n_1_67), .C1(n_31), .C2(n_1_66), .ZN(n_1_50));
   INV_X1 i_1_84 (.A(n_1_51), .ZN(n_16));
   AOI222_X1 i_1_85 (.A1(\temp1[12] [19]), .A2(n_1_68), .B1(\temp2[12] [19]), 
      .B2(n_1_67), .C1(n_32), .C2(n_1_66), .ZN(n_1_51));
   INV_X1 i_1_86 (.A(n_1_52), .ZN(n_17));
   AOI222_X1 i_1_87 (.A1(\temp1[12] [20]), .A2(n_1_68), .B1(\temp2[12] [20]), 
      .B2(n_1_67), .C1(n_33), .C2(n_1_66), .ZN(n_1_52));
   INV_X1 i_1_88 (.A(n_1_53), .ZN(n_18));
   AOI222_X1 i_1_89 (.A1(\temp1[12] [21]), .A2(n_1_68), .B1(\temp2[12] [21]), 
      .B2(n_1_67), .C1(n_34), .C2(n_1_66), .ZN(n_1_53));
   INV_X1 i_1_90 (.A(n_1_54), .ZN(n_19));
   AOI222_X1 i_1_91 (.A1(\temp1[12] [22]), .A2(n_1_68), .B1(\temp2[12] [22]), 
      .B2(n_1_67), .C1(n_35), .C2(n_1_66), .ZN(n_1_54));
   INV_X1 i_1_92 (.A(n_1_55), .ZN(n_20));
   AOI222_X1 i_1_93 (.A1(\temp1[12] [23]), .A2(n_1_68), .B1(\temp2[12] [23]), 
      .B2(n_1_67), .C1(n_36), .C2(n_1_66), .ZN(n_1_55));
   INV_X1 i_1_94 (.A(n_1_56), .ZN(n_21));
   AOI222_X1 i_1_95 (.A1(\temp1[12] [24]), .A2(n_1_68), .B1(\temp2[12] [24]), 
      .B2(n_1_67), .C1(n_37), .C2(n_1_66), .ZN(n_1_56));
   INV_X1 i_1_96 (.A(n_1_57), .ZN(n_22));
   AOI222_X1 i_1_97 (.A1(\temp1[12] [25]), .A2(n_1_68), .B1(\temp2[12] [25]), 
      .B2(n_1_67), .C1(n_38), .C2(n_1_66), .ZN(n_1_57));
   INV_X1 i_1_98 (.A(n_1_58), .ZN(n_23));
   AOI222_X1 i_1_99 (.A1(\temp1[12] [26]), .A2(n_1_68), .B1(\temp2[12] [26]), 
      .B2(n_1_67), .C1(n_39), .C2(n_1_66), .ZN(n_1_58));
   INV_X1 i_1_100 (.A(n_1_59), .ZN(n_24));
   AOI222_X1 i_1_101 (.A1(\temp1[12] [27]), .A2(n_1_68), .B1(\temp2[12] [27]), 
      .B2(n_1_67), .C1(n_40), .C2(n_1_66), .ZN(n_1_59));
   INV_X1 i_1_102 (.A(n_1_60), .ZN(n_25));
   AOI222_X1 i_1_103 (.A1(\temp1[12] [28]), .A2(n_1_68), .B1(\temp2[12] [28]), 
      .B2(n_1_67), .C1(n_41), .C2(n_1_66), .ZN(n_1_60));
   INV_X1 i_1_104 (.A(n_1_61), .ZN(n_26));
   AOI222_X1 i_1_105 (.A1(\temp1[12] [29]), .A2(n_1_68), .B1(\temp2[12] [29]), 
      .B2(n_1_67), .C1(n_42), .C2(n_1_66), .ZN(n_1_61));
   INV_X1 i_1_106 (.A(n_1_62), .ZN(n_27));
   AOI222_X1 i_1_107 (.A1(\temp1[12] [30]), .A2(n_1_68), .B1(\temp2[12] [30]), 
      .B2(n_1_67), .C1(n_43), .C2(n_1_66), .ZN(n_1_62));
   INV_X1 i_1_108 (.A(n_1_63), .ZN(n_28));
   AOI221_X1 i_1_109 (.A(n_1_65), .B1(\temp1[12] [31]), .B2(n_1_68), .C1(
      \temp2[12] [31]), .C2(n_1_67), .ZN(n_1_63));
   INV_X1 i_1_110 (.A(n_1_64), .ZN(n_29));
   AOI221_X1 i_1_111 (.A(n_1_65), .B1(\temp1[12] [32]), .B2(n_1_68), .C1(
      \temp2[12] [32]), .C2(n_1_67), .ZN(n_1_64));
   AND2_X1 i_1_112 (.A1(n_44), .A2(n_1_66), .ZN(n_1_65));
   NOR2_X1 i_1_113 (.A1(n_1_68), .A2(n_1_67), .ZN(n_1_66));
   NOR2_X1 i_1_114 (.A1(n_1_26), .A2(r[11]), .ZN(n_1_67));
   NOR2_X1 i_1_115 (.A1(r[12]), .A2(n_1_25), .ZN(n_1_68));
   INV_X1 i_1_116 (.A(n_1_69), .ZN(n_30));
   AOI222_X1 i_1_117 (.A1(\temp1[11] [18]), .A2(n_1_87), .B1(\temp2[11] [18]), 
      .B2(n_1_86), .C1(n_46), .C2(n_1_85), .ZN(n_1_69));
   INV_X1 i_1_118 (.A(n_1_70), .ZN(n_31));
   AOI222_X1 i_1_119 (.A1(\temp1[11] [19]), .A2(n_1_87), .B1(\temp2[11] [19]), 
      .B2(n_1_86), .C1(n_47), .C2(n_1_85), .ZN(n_1_70));
   INV_X1 i_1_120 (.A(n_1_71), .ZN(n_32));
   AOI222_X1 i_1_121 (.A1(\temp1[11] [20]), .A2(n_1_87), .B1(\temp2[11] [20]), 
      .B2(n_1_86), .C1(n_48), .C2(n_1_85), .ZN(n_1_71));
   INV_X1 i_1_122 (.A(n_1_72), .ZN(n_33));
   AOI222_X1 i_1_123 (.A1(\temp1[11] [21]), .A2(n_1_87), .B1(\temp2[11] [21]), 
      .B2(n_1_86), .C1(n_49), .C2(n_1_85), .ZN(n_1_72));
   INV_X1 i_1_124 (.A(n_1_73), .ZN(n_34));
   AOI222_X1 i_1_125 (.A1(\temp1[11] [22]), .A2(n_1_87), .B1(\temp2[11] [22]), 
      .B2(n_1_86), .C1(n_50), .C2(n_1_85), .ZN(n_1_73));
   INV_X1 i_1_126 (.A(n_1_74), .ZN(n_35));
   AOI222_X1 i_1_127 (.A1(\temp1[11] [23]), .A2(n_1_87), .B1(\temp2[11] [23]), 
      .B2(n_1_86), .C1(n_51), .C2(n_1_85), .ZN(n_1_74));
   INV_X1 i_1_128 (.A(n_1_75), .ZN(n_36));
   AOI222_X1 i_1_129 (.A1(\temp1[11] [24]), .A2(n_1_87), .B1(\temp2[11] [24]), 
      .B2(n_1_86), .C1(n_52), .C2(n_1_85), .ZN(n_1_75));
   INV_X1 i_1_130 (.A(n_1_76), .ZN(n_37));
   AOI222_X1 i_1_131 (.A1(\temp1[11] [25]), .A2(n_1_87), .B1(\temp2[11] [25]), 
      .B2(n_1_86), .C1(n_53), .C2(n_1_85), .ZN(n_1_76));
   INV_X1 i_1_132 (.A(n_1_77), .ZN(n_38));
   AOI222_X1 i_1_133 (.A1(\temp1[11] [26]), .A2(n_1_87), .B1(\temp2[11] [26]), 
      .B2(n_1_86), .C1(n_54), .C2(n_1_85), .ZN(n_1_77));
   INV_X1 i_1_134 (.A(n_1_78), .ZN(n_39));
   AOI222_X1 i_1_135 (.A1(\temp1[11] [27]), .A2(n_1_87), .B1(\temp2[11] [27]), 
      .B2(n_1_86), .C1(n_55), .C2(n_1_85), .ZN(n_1_78));
   INV_X1 i_1_136 (.A(n_1_79), .ZN(n_40));
   AOI222_X1 i_1_137 (.A1(\temp2[11] [28]), .A2(n_1_86), .B1(\temp1[11] [28]), 
      .B2(n_1_87), .C1(n_56), .C2(n_1_85), .ZN(n_1_79));
   INV_X1 i_1_138 (.A(n_1_80), .ZN(n_41));
   AOI222_X1 i_1_139 (.A1(\temp1[11] [29]), .A2(n_1_87), .B1(\temp2[11] [29]), 
      .B2(n_1_86), .C1(n_57), .C2(n_1_85), .ZN(n_1_80));
   INV_X1 i_1_140 (.A(n_1_81), .ZN(n_42));
   AOI222_X1 i_1_141 (.A1(\temp1[11] [30]), .A2(n_1_87), .B1(\temp2[11] [30]), 
      .B2(n_1_86), .C1(n_58), .C2(n_1_85), .ZN(n_1_81));
   INV_X1 i_1_142 (.A(n_1_82), .ZN(n_43));
   AOI221_X1 i_1_143 (.A(n_1_84), .B1(\temp1[11] [31]), .B2(n_1_87), .C1(
      \temp2[11] [31]), .C2(n_1_86), .ZN(n_1_82));
   INV_X1 i_1_144 (.A(n_1_83), .ZN(n_44));
   AOI221_X1 i_1_145 (.A(n_1_84), .B1(\temp1[11] [32]), .B2(n_1_87), .C1(
      \temp2[11] [32]), .C2(n_1_86), .ZN(n_1_83));
   AND2_X1 i_1_146 (.A1(n_59), .A2(n_1_85), .ZN(n_1_84));
   NOR2_X1 i_1_147 (.A1(n_1_87), .A2(n_1_86), .ZN(n_1_85));
   NOR2_X1 i_1_148 (.A1(n_1_25), .A2(r[10]), .ZN(n_1_86));
   NOR2_X1 i_1_149 (.A1(r[11]), .A2(n_1_24), .ZN(n_1_87));
   INV_X1 i_1_150 (.A(n_1_88), .ZN(n_45));
   AOI222_X1 i_1_151 (.A1(\temp2[10] [18]), .A2(n_1_105), .B1(\temp1[10] [18]), 
      .B2(n_1_106), .C1(n_61), .C2(n_1_104), .ZN(n_1_88));
   INV_X1 i_1_152 (.A(n_1_89), .ZN(n_46));
   AOI222_X1 i_1_153 (.A1(\temp1[10] [19]), .A2(n_1_106), .B1(\temp2[10] [19]), 
      .B2(n_1_105), .C1(n_62), .C2(n_1_104), .ZN(n_1_89));
   INV_X1 i_1_154 (.A(n_1_90), .ZN(n_47));
   AOI222_X1 i_1_155 (.A1(\temp1[10] [20]), .A2(n_1_106), .B1(\temp2[10] [20]), 
      .B2(n_1_105), .C1(n_63), .C2(n_1_104), .ZN(n_1_90));
   INV_X1 i_1_156 (.A(n_1_91), .ZN(n_48));
   AOI222_X1 i_1_157 (.A1(\temp1[10] [21]), .A2(n_1_106), .B1(\temp2[10] [21]), 
      .B2(n_1_105), .C1(n_64), .C2(n_1_104), .ZN(n_1_91));
   INV_X1 i_1_158 (.A(n_1_92), .ZN(n_49));
   AOI222_X1 i_1_159 (.A1(\temp1[10] [22]), .A2(n_1_106), .B1(\temp2[10] [22]), 
      .B2(n_1_105), .C1(n_65), .C2(n_1_104), .ZN(n_1_92));
   INV_X1 i_1_160 (.A(n_1_93), .ZN(n_50));
   AOI222_X1 i_1_161 (.A1(\temp1[10] [23]), .A2(n_1_106), .B1(\temp2[10] [23]), 
      .B2(n_1_105), .C1(n_66), .C2(n_1_104), .ZN(n_1_93));
   INV_X1 i_1_162 (.A(n_1_94), .ZN(n_51));
   AOI222_X1 i_1_163 (.A1(\temp1[10] [24]), .A2(n_1_106), .B1(\temp2[10] [24]), 
      .B2(n_1_105), .C1(n_67), .C2(n_1_104), .ZN(n_1_94));
   INV_X1 i_1_164 (.A(n_1_95), .ZN(n_52));
   AOI222_X1 i_1_165 (.A1(\temp1[10] [25]), .A2(n_1_106), .B1(\temp2[10] [25]), 
      .B2(n_1_105), .C1(n_68), .C2(n_1_104), .ZN(n_1_95));
   INV_X1 i_1_166 (.A(n_1_96), .ZN(n_53));
   AOI222_X1 i_1_167 (.A1(\temp1[10] [26]), .A2(n_1_106), .B1(\temp2[10] [26]), 
      .B2(n_1_105), .C1(n_69), .C2(n_1_104), .ZN(n_1_96));
   INV_X1 i_1_168 (.A(n_1_97), .ZN(n_54));
   AOI222_X1 i_1_169 (.A1(\temp1[10] [27]), .A2(n_1_106), .B1(\temp2[10] [27]), 
      .B2(n_1_105), .C1(n_70), .C2(n_1_104), .ZN(n_1_97));
   INV_X1 i_1_170 (.A(n_1_98), .ZN(n_55));
   AOI222_X1 i_1_171 (.A1(\temp2[10] [28]), .A2(n_1_105), .B1(\temp1[10] [28]), 
      .B2(n_1_106), .C1(n_71), .C2(n_1_104), .ZN(n_1_98));
   INV_X1 i_1_172 (.A(n_1_99), .ZN(n_56));
   AOI222_X1 i_1_173 (.A1(\temp2[10] [29]), .A2(n_1_105), .B1(\temp1[10] [29]), 
      .B2(n_1_106), .C1(n_72), .C2(n_1_104), .ZN(n_1_99));
   INV_X1 i_1_174 (.A(n_1_100), .ZN(n_57));
   AOI222_X1 i_1_175 (.A1(\temp1[10] [30]), .A2(n_1_106), .B1(\temp2[10] [30]), 
      .B2(n_1_105), .C1(n_73), .C2(n_1_104), .ZN(n_1_100));
   INV_X1 i_1_176 (.A(n_1_101), .ZN(n_58));
   AOI221_X1 i_1_177 (.A(n_1_103), .B1(\temp1[10] [31]), .B2(n_1_106), .C1(
      \temp2[10] [31]), .C2(n_1_105), .ZN(n_1_101));
   INV_X1 i_1_178 (.A(n_1_102), .ZN(n_59));
   AOI221_X1 i_1_179 (.A(n_1_103), .B1(\temp1[10] [32]), .B2(n_1_106), .C1(
      \temp2[10] [32]), .C2(n_1_105), .ZN(n_1_102));
   AND2_X1 i_1_180 (.A1(n_74), .A2(n_1_104), .ZN(n_1_103));
   NOR2_X1 i_1_181 (.A1(n_1_106), .A2(n_1_105), .ZN(n_1_104));
   NOR2_X1 i_1_182 (.A1(n_1_24), .A2(r[9]), .ZN(n_1_105));
   NOR2_X1 i_1_183 (.A1(r[10]), .A2(n_1_23), .ZN(n_1_106));
   INV_X1 i_1_184 (.A(n_1_107), .ZN(n_60));
   AOI222_X1 i_1_185 (.A1(\temp2[9] [18]), .A2(n_1_124), .B1(\temp1[9] [18]), 
      .B2(n_1_125), .C1(n_76), .C2(n_1_123), .ZN(n_1_107));
   INV_X1 i_1_186 (.A(n_1_108), .ZN(n_61));
   AOI222_X1 i_1_187 (.A1(\temp2[9] [19]), .A2(n_1_124), .B1(\temp1[9] [19]), 
      .B2(n_1_125), .C1(n_77), .C2(n_1_123), .ZN(n_1_108));
   INV_X1 i_1_188 (.A(n_1_109), .ZN(n_62));
   AOI222_X1 i_1_189 (.A1(\temp2[9] [20]), .A2(n_1_124), .B1(\temp1[9] [20]), 
      .B2(n_1_125), .C1(n_78), .C2(n_1_123), .ZN(n_1_109));
   INV_X1 i_1_190 (.A(n_1_110), .ZN(n_63));
   AOI222_X1 i_1_191 (.A1(\temp1[9] [21]), .A2(n_1_125), .B1(\temp2[9] [21]), 
      .B2(n_1_124), .C1(n_79), .C2(n_1_123), .ZN(n_1_110));
   INV_X1 i_1_192 (.A(n_1_111), .ZN(n_64));
   AOI222_X1 i_1_193 (.A1(\temp1[9] [22]), .A2(n_1_125), .B1(\temp2[9] [22]), 
      .B2(n_1_124), .C1(n_80), .C2(n_1_123), .ZN(n_1_111));
   INV_X1 i_1_194 (.A(n_1_112), .ZN(n_65));
   AOI222_X1 i_1_195 (.A1(\temp1[9] [23]), .A2(n_1_125), .B1(\temp2[9] [23]), 
      .B2(n_1_124), .C1(n_81), .C2(n_1_123), .ZN(n_1_112));
   INV_X1 i_1_196 (.A(n_1_113), .ZN(n_66));
   AOI222_X1 i_1_197 (.A1(\temp1[9] [24]), .A2(n_1_125), .B1(\temp2[9] [24]), 
      .B2(n_1_124), .C1(n_82), .C2(n_1_123), .ZN(n_1_113));
   INV_X1 i_1_198 (.A(n_1_114), .ZN(n_67));
   AOI222_X1 i_1_199 (.A1(\temp1[9] [25]), .A2(n_1_125), .B1(\temp2[9] [25]), 
      .B2(n_1_124), .C1(n_83), .C2(n_1_123), .ZN(n_1_114));
   INV_X1 i_1_200 (.A(n_1_115), .ZN(n_68));
   AOI222_X1 i_1_201 (.A1(\temp1[9] [26]), .A2(n_1_125), .B1(\temp2[9] [26]), 
      .B2(n_1_124), .C1(n_84), .C2(n_1_123), .ZN(n_1_115));
   INV_X1 i_1_202 (.A(n_1_116), .ZN(n_69));
   AOI222_X1 i_1_203 (.A1(\temp1[9] [27]), .A2(n_1_125), .B1(\temp2[9] [27]), 
      .B2(n_1_124), .C1(n_85), .C2(n_1_123), .ZN(n_1_116));
   INV_X1 i_1_204 (.A(n_1_117), .ZN(n_70));
   AOI222_X1 i_1_205 (.A1(\temp2[9] [28]), .A2(n_1_124), .B1(\temp1[9] [28]), 
      .B2(n_1_125), .C1(n_86), .C2(n_1_123), .ZN(n_1_117));
   INV_X1 i_1_206 (.A(n_1_118), .ZN(n_71));
   AOI222_X1 i_1_207 (.A1(\temp2[9] [29]), .A2(n_1_124), .B1(\temp1[9] [29]), 
      .B2(n_1_125), .C1(n_87), .C2(n_1_123), .ZN(n_1_118));
   INV_X1 i_1_208 (.A(n_1_119), .ZN(n_72));
   AOI222_X1 i_1_209 (.A1(\temp2[9] [30]), .A2(n_1_124), .B1(\temp1[9] [30]), 
      .B2(n_1_125), .C1(n_88), .C2(n_1_123), .ZN(n_1_119));
   INV_X1 i_1_210 (.A(n_1_120), .ZN(n_73));
   AOI221_X1 i_1_211 (.A(n_1_122), .B1(\temp1[9] [31]), .B2(n_1_125), .C1(
      \temp2[9] [31]), .C2(n_1_124), .ZN(n_1_120));
   INV_X1 i_1_212 (.A(n_1_121), .ZN(n_74));
   AOI221_X1 i_1_213 (.A(n_1_122), .B1(\temp1[9] [32]), .B2(n_1_125), .C1(
      \temp2[9] [32]), .C2(n_1_124), .ZN(n_1_121));
   AND2_X1 i_1_214 (.A1(n_89), .A2(n_1_123), .ZN(n_1_122));
   NOR2_X1 i_1_215 (.A1(n_1_125), .A2(n_1_124), .ZN(n_1_123));
   NOR2_X1 i_1_216 (.A1(n_1_23), .A2(r[8]), .ZN(n_1_124));
   NOR2_X1 i_1_217 (.A1(r[9]), .A2(n_1_22), .ZN(n_1_125));
   INV_X1 i_1_218 (.A(n_1_126), .ZN(n_75));
   AOI222_X1 i_1_219 (.A1(\temp2[8] [18]), .A2(n_1_143), .B1(\temp1[8] [18]), 
      .B2(n_1_144), .C1(n_91), .C2(n_1_142), .ZN(n_1_126));
   INV_X1 i_1_220 (.A(n_1_127), .ZN(n_76));
   AOI222_X1 i_1_221 (.A1(\temp2[8] [19]), .A2(n_1_143), .B1(\temp1[8] [19]), 
      .B2(n_1_144), .C1(n_92), .C2(n_1_142), .ZN(n_1_127));
   INV_X1 i_1_222 (.A(n_1_128), .ZN(n_77));
   AOI222_X1 i_1_223 (.A1(\temp2[8] [20]), .A2(n_1_143), .B1(\temp1[8] [20]), 
      .B2(n_1_144), .C1(n_93), .C2(n_1_142), .ZN(n_1_128));
   INV_X1 i_1_224 (.A(n_1_129), .ZN(n_78));
   AOI222_X1 i_1_225 (.A1(\temp2[8] [21]), .A2(n_1_143), .B1(\temp1[8] [21]), 
      .B2(n_1_144), .C1(n_94), .C2(n_1_142), .ZN(n_1_129));
   INV_X1 i_1_226 (.A(n_1_130), .ZN(n_79));
   AOI222_X1 i_1_227 (.A1(\temp1[8] [22]), .A2(n_1_144), .B1(\temp2[8] [22]), 
      .B2(n_1_143), .C1(n_95), .C2(n_1_142), .ZN(n_1_130));
   INV_X1 i_1_228 (.A(n_1_131), .ZN(n_80));
   AOI222_X1 i_1_229 (.A1(\temp1[8] [23]), .A2(n_1_144), .B1(\temp2[8] [23]), 
      .B2(n_1_143), .C1(n_96), .C2(n_1_142), .ZN(n_1_131));
   INV_X1 i_1_230 (.A(n_1_132), .ZN(n_81));
   AOI222_X1 i_1_231 (.A1(\temp1[8] [24]), .A2(n_1_144), .B1(\temp2[8] [24]), 
      .B2(n_1_143), .C1(n_97), .C2(n_1_142), .ZN(n_1_132));
   INV_X1 i_1_232 (.A(n_1_133), .ZN(n_82));
   AOI222_X1 i_1_233 (.A1(\temp1[8] [25]), .A2(n_1_144), .B1(\temp2[8] [25]), 
      .B2(n_1_143), .C1(n_98), .C2(n_1_142), .ZN(n_1_133));
   INV_X1 i_1_234 (.A(n_1_134), .ZN(n_83));
   AOI222_X1 i_1_235 (.A1(\temp1[8] [26]), .A2(n_1_144), .B1(\temp2[8] [26]), 
      .B2(n_1_143), .C1(n_99), .C2(n_1_142), .ZN(n_1_134));
   INV_X1 i_1_236 (.A(n_1_135), .ZN(n_84));
   AOI222_X1 i_1_237 (.A1(\temp1[8] [27]), .A2(n_1_144), .B1(\temp2[8] [27]), 
      .B2(n_1_143), .C1(n_100), .C2(n_1_142), .ZN(n_1_135));
   INV_X1 i_1_238 (.A(n_1_136), .ZN(n_85));
   AOI222_X1 i_1_239 (.A1(\temp2[8] [28]), .A2(n_1_143), .B1(\temp1[8] [28]), 
      .B2(n_1_144), .C1(n_101), .C2(n_1_142), .ZN(n_1_136));
   INV_X1 i_1_240 (.A(n_1_137), .ZN(n_86));
   AOI222_X1 i_1_241 (.A1(\temp2[8] [29]), .A2(n_1_143), .B1(\temp1[8] [29]), 
      .B2(n_1_144), .C1(n_102), .C2(n_1_142), .ZN(n_1_137));
   INV_X1 i_1_242 (.A(n_1_138), .ZN(n_87));
   AOI222_X1 i_1_243 (.A1(\temp2[8] [30]), .A2(n_1_143), .B1(\temp1[8] [30]), 
      .B2(n_1_144), .C1(n_103), .C2(n_1_142), .ZN(n_1_138));
   INV_X1 i_1_244 (.A(n_1_139), .ZN(n_88));
   AOI221_X1 i_1_245 (.A(n_1_141), .B1(\temp1[8] [31]), .B2(n_1_144), .C1(
      \temp2[8] [31]), .C2(n_1_143), .ZN(n_1_139));
   INV_X1 i_1_246 (.A(n_1_140), .ZN(n_89));
   AOI221_X1 i_1_247 (.A(n_1_141), .B1(\temp1[8] [32]), .B2(n_1_144), .C1(
      \temp2[8] [32]), .C2(n_1_143), .ZN(n_1_140));
   AND2_X1 i_1_248 (.A1(n_104), .A2(n_1_142), .ZN(n_1_141));
   NOR2_X1 i_1_249 (.A1(n_1_144), .A2(n_1_143), .ZN(n_1_142));
   NOR2_X1 i_1_250 (.A1(n_1_22), .A2(r[7]), .ZN(n_1_143));
   NOR2_X1 i_1_251 (.A1(r[8]), .A2(n_1_21), .ZN(n_1_144));
   INV_X1 i_1_252 (.A(n_1_145), .ZN(n_90));
   AOI222_X1 i_1_253 (.A1(\temp2[7] [18]), .A2(n_1_162), .B1(\temp1[7] [18]), 
      .B2(n_1_163), .C1(n_106), .C2(n_1_161), .ZN(n_1_145));
   INV_X1 i_1_254 (.A(n_1_146), .ZN(n_91));
   AOI222_X1 i_1_255 (.A1(\temp2[7] [19]), .A2(n_1_162), .B1(\temp1[7] [19]), 
      .B2(n_1_163), .C1(n_107), .C2(n_1_161), .ZN(n_1_146));
   INV_X1 i_1_256 (.A(n_1_147), .ZN(n_92));
   AOI222_X1 i_1_257 (.A1(\temp2[7] [20]), .A2(n_1_162), .B1(\temp1[7] [20]), 
      .B2(n_1_163), .C1(n_108), .C2(n_1_161), .ZN(n_1_147));
   INV_X1 i_1_258 (.A(n_1_148), .ZN(n_93));
   AOI222_X1 i_1_259 (.A1(\temp2[7] [21]), .A2(n_1_162), .B1(\temp1[7] [21]), 
      .B2(n_1_163), .C1(n_109), .C2(n_1_161), .ZN(n_1_148));
   INV_X1 i_1_260 (.A(n_1_149), .ZN(n_94));
   AOI222_X1 i_1_261 (.A1(\temp2[7] [22]), .A2(n_1_162), .B1(\temp1[7] [22]), 
      .B2(n_1_163), .C1(n_110), .C2(n_1_161), .ZN(n_1_149));
   INV_X1 i_1_262 (.A(n_1_150), .ZN(n_95));
   AOI222_X1 i_1_263 (.A1(\temp2[7] [23]), .A2(n_1_162), .B1(\temp1[7] [23]), 
      .B2(n_1_163), .C1(n_111), .C2(n_1_161), .ZN(n_1_150));
   INV_X1 i_1_264 (.A(n_1_151), .ZN(n_96));
   AOI222_X1 i_1_265 (.A1(\temp1[7] [24]), .A2(n_1_163), .B1(\temp2[7] [24]), 
      .B2(n_1_162), .C1(n_112), .C2(n_1_161), .ZN(n_1_151));
   INV_X1 i_1_266 (.A(n_1_152), .ZN(n_97));
   AOI222_X1 i_1_267 (.A1(\temp1[7] [25]), .A2(n_1_163), .B1(\temp2[7] [25]), 
      .B2(n_1_162), .C1(n_113), .C2(n_1_161), .ZN(n_1_152));
   INV_X1 i_1_268 (.A(n_1_153), .ZN(n_98));
   AOI222_X1 i_1_269 (.A1(\temp1[7] [26]), .A2(n_1_163), .B1(\temp2[7] [26]), 
      .B2(n_1_162), .C1(n_114), .C2(n_1_161), .ZN(n_1_153));
   INV_X1 i_1_270 (.A(n_1_154), .ZN(n_99));
   AOI222_X1 i_1_271 (.A1(\temp1[7] [27]), .A2(n_1_163), .B1(\temp2[7] [27]), 
      .B2(n_1_162), .C1(n_115), .C2(n_1_161), .ZN(n_1_154));
   INV_X1 i_1_272 (.A(n_1_155), .ZN(n_100));
   AOI222_X1 i_1_273 (.A1(\temp2[7] [28]), .A2(n_1_162), .B1(\temp1[7] [28]), 
      .B2(n_1_163), .C1(n_116), .C2(n_1_161), .ZN(n_1_155));
   INV_X1 i_1_274 (.A(n_1_156), .ZN(n_101));
   AOI222_X1 i_1_275 (.A1(\temp2[7] [29]), .A2(n_1_162), .B1(\temp1[7] [29]), 
      .B2(n_1_163), .C1(n_117), .C2(n_1_161), .ZN(n_1_156));
   INV_X1 i_1_276 (.A(n_1_157), .ZN(n_102));
   AOI222_X1 i_1_277 (.A1(\temp2[7] [30]), .A2(n_1_162), .B1(\temp1[7] [30]), 
      .B2(n_1_163), .C1(n_118), .C2(n_1_161), .ZN(n_1_157));
   INV_X1 i_1_278 (.A(n_1_158), .ZN(n_103));
   AOI221_X1 i_1_279 (.A(n_1_160), .B1(\temp1[7] [31]), .B2(n_1_163), .C1(
      \temp2[7] [31]), .C2(n_1_162), .ZN(n_1_158));
   INV_X1 i_1_280 (.A(n_1_159), .ZN(n_104));
   AOI221_X1 i_1_281 (.A(n_1_160), .B1(\temp1[7] [32]), .B2(n_1_163), .C1(
      \temp2[7] [32]), .C2(n_1_162), .ZN(n_1_159));
   AND2_X1 i_1_282 (.A1(n_119), .A2(n_1_161), .ZN(n_1_160));
   NOR2_X1 i_1_283 (.A1(n_1_163), .A2(n_1_162), .ZN(n_1_161));
   NOR2_X1 i_1_284 (.A1(n_1_21), .A2(r[6]), .ZN(n_1_162));
   NOR2_X1 i_1_285 (.A1(r[7]), .A2(n_1_20), .ZN(n_1_163));
   INV_X1 i_1_286 (.A(n_1_164), .ZN(n_105));
   AOI222_X1 i_1_287 (.A1(\temp2[6] [18]), .A2(n_1_181), .B1(\temp1[6] [18]), 
      .B2(n_1_182), .C1(n_121), .C2(n_1_180), .ZN(n_1_164));
   INV_X1 i_1_288 (.A(n_1_165), .ZN(n_106));
   AOI222_X1 i_1_289 (.A1(\temp2[6] [19]), .A2(n_1_181), .B1(\temp1[6] [19]), 
      .B2(n_1_182), .C1(n_122), .C2(n_1_180), .ZN(n_1_165));
   INV_X1 i_1_290 (.A(n_1_166), .ZN(n_107));
   AOI222_X1 i_1_291 (.A1(\temp2[6] [20]), .A2(n_1_181), .B1(\temp1[6] [20]), 
      .B2(n_1_182), .C1(n_123), .C2(n_1_180), .ZN(n_1_166));
   INV_X1 i_1_292 (.A(n_1_167), .ZN(n_108));
   AOI222_X1 i_1_293 (.A1(\temp2[6] [21]), .A2(n_1_181), .B1(\temp1[6] [21]), 
      .B2(n_1_182), .C1(n_124), .C2(n_1_180), .ZN(n_1_167));
   INV_X1 i_1_294 (.A(n_1_168), .ZN(n_109));
   AOI222_X1 i_1_295 (.A1(\temp2[6] [22]), .A2(n_1_181), .B1(\temp1[6] [22]), 
      .B2(n_1_182), .C1(n_125), .C2(n_1_180), .ZN(n_1_168));
   INV_X1 i_1_296 (.A(n_1_169), .ZN(n_110));
   AOI222_X1 i_1_297 (.A1(\temp2[6] [23]), .A2(n_1_181), .B1(\temp1[6] [23]), 
      .B2(n_1_182), .C1(n_126), .C2(n_1_180), .ZN(n_1_169));
   INV_X1 i_1_298 (.A(n_1_170), .ZN(n_111));
   AOI222_X1 i_1_299 (.A1(\temp2[6] [24]), .A2(n_1_181), .B1(\temp1[6] [24]), 
      .B2(n_1_182), .C1(n_127), .C2(n_1_180), .ZN(n_1_170));
   INV_X1 i_1_300 (.A(n_1_171), .ZN(n_112));
   AOI222_X1 i_1_301 (.A1(\temp1[6] [25]), .A2(n_1_182), .B1(\temp2[6] [25]), 
      .B2(n_1_181), .C1(n_128), .C2(n_1_180), .ZN(n_1_171));
   INV_X1 i_1_302 (.A(n_1_172), .ZN(n_113));
   AOI222_X1 i_1_303 (.A1(\temp1[6] [26]), .A2(n_1_182), .B1(\temp2[6] [26]), 
      .B2(n_1_181), .C1(n_129), .C2(n_1_180), .ZN(n_1_172));
   INV_X1 i_1_304 (.A(n_1_173), .ZN(n_114));
   AOI222_X1 i_1_305 (.A1(\temp1[6] [27]), .A2(n_1_182), .B1(\temp2[6] [27]), 
      .B2(n_1_181), .C1(n_130), .C2(n_1_180), .ZN(n_1_173));
   INV_X1 i_1_306 (.A(n_1_174), .ZN(n_115));
   AOI222_X1 i_1_307 (.A1(\temp2[6] [28]), .A2(n_1_181), .B1(\temp1[6] [28]), 
      .B2(n_1_182), .C1(n_131), .C2(n_1_180), .ZN(n_1_174));
   INV_X1 i_1_308 (.A(n_1_175), .ZN(n_116));
   AOI222_X1 i_1_309 (.A1(\temp2[6] [29]), .A2(n_1_181), .B1(\temp1[6] [29]), 
      .B2(n_1_182), .C1(n_132), .C2(n_1_180), .ZN(n_1_175));
   INV_X1 i_1_310 (.A(n_1_176), .ZN(n_117));
   AOI222_X1 i_1_311 (.A1(\temp2[6] [30]), .A2(n_1_181), .B1(\temp1[6] [30]), 
      .B2(n_1_182), .C1(n_133), .C2(n_1_180), .ZN(n_1_176));
   INV_X1 i_1_312 (.A(n_1_177), .ZN(n_118));
   AOI221_X1 i_1_313 (.A(n_1_179), .B1(\temp1[6] [31]), .B2(n_1_182), .C1(
      \temp2[6] [31]), .C2(n_1_181), .ZN(n_1_177));
   INV_X1 i_1_314 (.A(n_1_178), .ZN(n_119));
   AOI221_X1 i_1_315 (.A(n_1_179), .B1(\temp1[6] [32]), .B2(n_1_182), .C1(
      \temp2[6] [32]), .C2(n_1_181), .ZN(n_1_178));
   AND2_X1 i_1_316 (.A1(n_134), .A2(n_1_180), .ZN(n_1_179));
   NOR2_X1 i_1_317 (.A1(n_1_182), .A2(n_1_181), .ZN(n_1_180));
   NOR2_X1 i_1_318 (.A1(n_1_20), .A2(r[5]), .ZN(n_1_181));
   NOR2_X1 i_1_319 (.A1(r[6]), .A2(n_1_19), .ZN(n_1_182));
   INV_X1 i_1_320 (.A(n_1_183), .ZN(n_120));
   AOI222_X1 i_1_321 (.A1(\temp2[5] [18]), .A2(n_1_200), .B1(\temp1[5] [18]), 
      .B2(n_1_201), .C1(n_136), .C2(n_1_199), .ZN(n_1_183));
   INV_X1 i_1_322 (.A(n_1_184), .ZN(n_121));
   AOI222_X1 i_1_323 (.A1(\temp2[5] [19]), .A2(n_1_200), .B1(\temp1[5] [19]), 
      .B2(n_1_201), .C1(n_137), .C2(n_1_199), .ZN(n_1_184));
   INV_X1 i_1_324 (.A(n_1_185), .ZN(n_122));
   AOI222_X1 i_1_325 (.A1(\temp2[5] [20]), .A2(n_1_200), .B1(\temp1[5] [20]), 
      .B2(n_1_201), .C1(n_138), .C2(n_1_199), .ZN(n_1_185));
   INV_X1 i_1_326 (.A(n_1_186), .ZN(n_123));
   AOI222_X1 i_1_327 (.A1(\temp2[5] [21]), .A2(n_1_200), .B1(\temp1[5] [21]), 
      .B2(n_1_201), .C1(n_139), .C2(n_1_199), .ZN(n_1_186));
   INV_X1 i_1_328 (.A(n_1_187), .ZN(n_124));
   AOI222_X1 i_1_329 (.A1(\temp2[5] [22]), .A2(n_1_200), .B1(\temp1[5] [22]), 
      .B2(n_1_201), .C1(n_140), .C2(n_1_199), .ZN(n_1_187));
   INV_X1 i_1_330 (.A(n_1_188), .ZN(n_125));
   AOI222_X1 i_1_331 (.A1(\temp2[5] [23]), .A2(n_1_200), .B1(\temp1[5] [23]), 
      .B2(n_1_201), .C1(n_141), .C2(n_1_199), .ZN(n_1_188));
   INV_X1 i_1_332 (.A(n_1_189), .ZN(n_126));
   AOI222_X1 i_1_333 (.A1(\temp2[5] [24]), .A2(n_1_200), .B1(\temp1[5] [24]), 
      .B2(n_1_201), .C1(n_142), .C2(n_1_199), .ZN(n_1_189));
   INV_X1 i_1_334 (.A(n_1_190), .ZN(n_127));
   AOI222_X1 i_1_335 (.A1(\temp2[5] [25]), .A2(n_1_200), .B1(\temp1[5] [25]), 
      .B2(n_1_201), .C1(n_143), .C2(n_1_199), .ZN(n_1_190));
   INV_X1 i_1_336 (.A(n_1_191), .ZN(n_128));
   AOI222_X1 i_1_337 (.A1(\temp2[5] [26]), .A2(n_1_200), .B1(\temp1[5] [26]), 
      .B2(n_1_201), .C1(n_144), .C2(n_1_199), .ZN(n_1_191));
   INV_X1 i_1_338 (.A(n_1_192), .ZN(n_129));
   AOI222_X1 i_1_339 (.A1(\temp2[5] [27]), .A2(n_1_200), .B1(\temp1[5] [27]), 
      .B2(n_1_201), .C1(n_145), .C2(n_1_199), .ZN(n_1_192));
   INV_X1 i_1_340 (.A(n_1_193), .ZN(n_130));
   AOI222_X1 i_1_341 (.A1(\temp2[5] [28]), .A2(n_1_200), .B1(\temp1[5] [28]), 
      .B2(n_1_201), .C1(n_146), .C2(n_1_199), .ZN(n_1_193));
   INV_X1 i_1_342 (.A(n_1_194), .ZN(n_131));
   AOI222_X1 i_1_343 (.A1(\temp2[5] [29]), .A2(n_1_200), .B1(\temp1[5] [29]), 
      .B2(n_1_201), .C1(n_147), .C2(n_1_199), .ZN(n_1_194));
   INV_X1 i_1_344 (.A(n_1_195), .ZN(n_132));
   AOI222_X1 i_1_345 (.A1(\temp2[5] [30]), .A2(n_1_200), .B1(\temp1[5] [30]), 
      .B2(n_1_201), .C1(n_148), .C2(n_1_199), .ZN(n_1_195));
   INV_X1 i_1_346 (.A(n_1_196), .ZN(n_133));
   AOI221_X1 i_1_347 (.A(n_1_198), .B1(\temp1[5] [31]), .B2(n_1_201), .C1(
      \temp2[5] [31]), .C2(n_1_200), .ZN(n_1_196));
   INV_X1 i_1_348 (.A(n_1_197), .ZN(n_134));
   AOI221_X1 i_1_349 (.A(n_1_198), .B1(\temp1[5] [32]), .B2(n_1_201), .C1(
      \temp2[5] [32]), .C2(n_1_200), .ZN(n_1_197));
   AND2_X1 i_1_350 (.A1(n_149), .A2(n_1_199), .ZN(n_1_198));
   NOR2_X1 i_1_351 (.A1(n_1_201), .A2(n_1_200), .ZN(n_1_199));
   NOR2_X1 i_1_352 (.A1(n_1_19), .A2(r[4]), .ZN(n_1_200));
   NOR2_X1 i_1_353 (.A1(r[5]), .A2(n_1_18), .ZN(n_1_201));
   INV_X1 i_1_354 (.A(n_1_202), .ZN(n_135));
   AOI222_X1 i_1_355 (.A1(\temp2[4] [18]), .A2(n_1_219), .B1(\temp1[4] [18]), 
      .B2(n_1_220), .C1(n_151), .C2(n_1_218), .ZN(n_1_202));
   INV_X1 i_1_356 (.A(n_1_203), .ZN(n_136));
   AOI222_X1 i_1_357 (.A1(\temp2[4] [19]), .A2(n_1_219), .B1(\temp1[4] [19]), 
      .B2(n_1_220), .C1(n_152), .C2(n_1_218), .ZN(n_1_203));
   INV_X1 i_1_358 (.A(n_1_204), .ZN(n_137));
   AOI222_X1 i_1_359 (.A1(\temp1[4] [20]), .A2(n_1_220), .B1(\temp2[4] [20]), 
      .B2(n_1_219), .C1(n_153), .C2(n_1_218), .ZN(n_1_204));
   INV_X1 i_1_360 (.A(n_1_205), .ZN(n_138));
   AOI222_X1 i_1_361 (.A1(\temp1[4] [21]), .A2(n_1_220), .B1(\temp2[4] [21]), 
      .B2(n_1_219), .C1(n_154), .C2(n_1_218), .ZN(n_1_205));
   INV_X1 i_1_362 (.A(n_1_206), .ZN(n_139));
   AOI222_X1 i_1_363 (.A1(\temp1[4] [22]), .A2(n_1_220), .B1(\temp2[4] [22]), 
      .B2(n_1_219), .C1(n_155), .C2(n_1_218), .ZN(n_1_206));
   INV_X1 i_1_364 (.A(n_1_207), .ZN(n_140));
   AOI222_X1 i_1_365 (.A1(\temp1[4] [23]), .A2(n_1_220), .B1(\temp2[4] [23]), 
      .B2(n_1_219), .C1(n_156), .C2(n_1_218), .ZN(n_1_207));
   INV_X1 i_1_366 (.A(n_1_208), .ZN(n_141));
   AOI222_X1 i_1_367 (.A1(\temp1[4] [24]), .A2(n_1_220), .B1(\temp2[4] [24]), 
      .B2(n_1_219), .C1(n_157), .C2(n_1_218), .ZN(n_1_208));
   INV_X1 i_1_368 (.A(n_1_209), .ZN(n_142));
   AOI222_X1 i_1_369 (.A1(\temp1[4] [25]), .A2(n_1_220), .B1(\temp2[4] [25]), 
      .B2(n_1_219), .C1(n_158), .C2(n_1_218), .ZN(n_1_209));
   INV_X1 i_1_370 (.A(n_1_210), .ZN(n_143));
   AOI222_X1 i_1_371 (.A1(\temp1[4] [26]), .A2(n_1_220), .B1(\temp2[4] [26]), 
      .B2(n_1_219), .C1(n_159), .C2(n_1_218), .ZN(n_1_210));
   INV_X1 i_1_372 (.A(n_1_211), .ZN(n_144));
   AOI222_X1 i_1_373 (.A1(\temp1[4] [27]), .A2(n_1_220), .B1(\temp2[4] [27]), 
      .B2(n_1_219), .C1(n_160), .C2(n_1_218), .ZN(n_1_211));
   INV_X1 i_1_374 (.A(n_1_212), .ZN(n_145));
   AOI222_X1 i_1_375 (.A1(\temp1[4] [28]), .A2(n_1_220), .B1(\temp2[4] [28]), 
      .B2(n_1_219), .C1(n_161), .C2(n_1_218), .ZN(n_1_212));
   INV_X1 i_1_376 (.A(n_1_213), .ZN(n_146));
   AOI222_X1 i_1_377 (.A1(\temp2[4] [29]), .A2(n_1_219), .B1(\temp1[4] [29]), 
      .B2(n_1_220), .C1(n_162), .C2(n_1_218), .ZN(n_1_213));
   INV_X1 i_1_378 (.A(n_1_214), .ZN(n_147));
   AOI222_X1 i_1_379 (.A1(\temp2[4] [30]), .A2(n_1_219), .B1(\temp1[4] [30]), 
      .B2(n_1_220), .C1(n_163), .C2(n_1_218), .ZN(n_1_214));
   INV_X1 i_1_380 (.A(n_1_215), .ZN(n_148));
   AOI221_X1 i_1_381 (.A(n_1_217), .B1(\temp1[4] [31]), .B2(n_1_220), .C1(
      \temp2[4] [31]), .C2(n_1_219), .ZN(n_1_215));
   INV_X1 i_1_382 (.A(n_1_216), .ZN(n_149));
   AOI221_X1 i_1_383 (.A(n_1_217), .B1(\temp1[4] [32]), .B2(n_1_220), .C1(
      \temp2[4] [32]), .C2(n_1_219), .ZN(n_1_216));
   AND2_X1 i_1_384 (.A1(n_164), .A2(n_1_218), .ZN(n_1_217));
   NOR2_X1 i_1_385 (.A1(n_1_220), .A2(n_1_219), .ZN(n_1_218));
   NOR2_X1 i_1_386 (.A1(n_1_18), .A2(r[3]), .ZN(n_1_219));
   NOR2_X1 i_1_387 (.A1(r[4]), .A2(n_1_17), .ZN(n_1_220));
   INV_X1 i_1_388 (.A(n_1_221), .ZN(n_150));
   AOI222_X1 i_1_389 (.A1(\temp1[3] [18]), .A2(n_1_239), .B1(\temp2[3] [18]), 
      .B2(n_1_238), .C1(n_166), .C2(n_1_237), .ZN(n_1_221));
   INV_X1 i_1_390 (.A(n_1_222), .ZN(n_151));
   AOI222_X1 i_1_391 (.A1(\temp2[3] [19]), .A2(n_1_238), .B1(\temp1[3] [19]), 
      .B2(n_1_239), .C1(n_167), .C2(n_1_237), .ZN(n_1_222));
   INV_X1 i_1_392 (.A(n_1_223), .ZN(n_152));
   AOI222_X1 i_1_393 (.A1(\temp2[3] [20]), .A2(n_1_238), .B1(\temp1[3] [20]), 
      .B2(n_1_239), .C1(n_168), .C2(n_1_237), .ZN(n_1_223));
   INV_X1 i_1_394 (.A(n_1_224), .ZN(n_153));
   AOI222_X1 i_1_395 (.A1(\temp2[3] [21]), .A2(n_1_238), .B1(\temp1[3] [21]), 
      .B2(n_1_239), .C1(n_169), .C2(n_1_237), .ZN(n_1_224));
   INV_X1 i_1_396 (.A(n_1_225), .ZN(n_154));
   AOI222_X1 i_1_397 (.A1(\temp2[3] [22]), .A2(n_1_238), .B1(\temp1[3] [22]), 
      .B2(n_1_239), .C1(n_170), .C2(n_1_237), .ZN(n_1_225));
   INV_X1 i_1_398 (.A(n_1_226), .ZN(n_155));
   AOI222_X1 i_1_399 (.A1(\temp2[3] [23]), .A2(n_1_238), .B1(\temp1[3] [23]), 
      .B2(n_1_239), .C1(n_171), .C2(n_1_237), .ZN(n_1_226));
   INV_X1 i_1_400 (.A(n_1_227), .ZN(n_156));
   AOI222_X1 i_1_401 (.A1(\temp2[3] [24]), .A2(n_1_238), .B1(\temp1[3] [24]), 
      .B2(n_1_239), .C1(n_172), .C2(n_1_237), .ZN(n_1_227));
   INV_X1 i_1_402 (.A(n_1_228), .ZN(n_157));
   AOI222_X1 i_1_403 (.A1(\temp2[3] [25]), .A2(n_1_238), .B1(\temp1[3] [25]), 
      .B2(n_1_239), .C1(n_173), .C2(n_1_237), .ZN(n_1_228));
   INV_X1 i_1_404 (.A(n_1_229), .ZN(n_158));
   AOI222_X1 i_1_405 (.A1(\temp2[3] [26]), .A2(n_1_238), .B1(\temp1[3] [26]), 
      .B2(n_1_239), .C1(n_174), .C2(n_1_237), .ZN(n_1_229));
   INV_X1 i_1_406 (.A(n_1_230), .ZN(n_159));
   AOI222_X1 i_1_407 (.A1(\temp2[3] [27]), .A2(n_1_238), .B1(\temp1[3] [27]), 
      .B2(n_1_239), .C1(n_175), .C2(n_1_237), .ZN(n_1_230));
   INV_X1 i_1_408 (.A(n_1_231), .ZN(n_160));
   AOI222_X1 i_1_409 (.A1(\temp2[3] [28]), .A2(n_1_238), .B1(\temp1[3] [28]), 
      .B2(n_1_239), .C1(n_176), .C2(n_1_237), .ZN(n_1_231));
   INV_X1 i_1_410 (.A(n_1_232), .ZN(n_161));
   AOI222_X1 i_1_411 (.A1(\temp2[3] [29]), .A2(n_1_238), .B1(\temp1[3] [29]), 
      .B2(n_1_239), .C1(n_177), .C2(n_1_237), .ZN(n_1_232));
   INV_X1 i_1_412 (.A(n_1_233), .ZN(n_162));
   AOI222_X1 i_1_413 (.A1(\temp2[3] [30]), .A2(n_1_238), .B1(\temp1[3] [30]), 
      .B2(n_1_239), .C1(n_178), .C2(n_1_237), .ZN(n_1_233));
   INV_X1 i_1_414 (.A(n_1_234), .ZN(n_163));
   AOI221_X1 i_1_415 (.A(n_1_236), .B1(\temp1[3] [31]), .B2(n_1_239), .C1(
      \temp2[3] [31]), .C2(n_1_238), .ZN(n_1_234));
   INV_X1 i_1_416 (.A(n_1_235), .ZN(n_164));
   AOI221_X1 i_1_417 (.A(n_1_236), .B1(\temp1[3] [32]), .B2(n_1_239), .C1(
      \temp2[3] [32]), .C2(n_1_238), .ZN(n_1_235));
   AND2_X1 i_1_418 (.A1(n_179), .A2(n_1_237), .ZN(n_1_236));
   NOR2_X1 i_1_419 (.A1(n_1_239), .A2(n_1_238), .ZN(n_1_237));
   NOR2_X1 i_1_420 (.A1(n_1_17), .A2(r[2]), .ZN(n_1_238));
   NOR2_X1 i_1_421 (.A1(r[3]), .A2(n_1_16), .ZN(n_1_239));
   INV_X1 i_1_422 (.A(n_1_240), .ZN(n_165));
   AOI222_X1 i_1_423 (.A1(\temp2[2] [18]), .A2(n_1_257), .B1(\temp1[2] [18]), 
      .B2(n_1_258), .C1(n_181), .C2(n_1_256), .ZN(n_1_240));
   INV_X1 i_1_424 (.A(n_1_241), .ZN(n_166));
   AOI222_X1 i_1_425 (.A1(\temp2[2] [19]), .A2(n_1_257), .B1(\temp1[2] [19]), 
      .B2(n_1_258), .C1(n_182), .C2(n_1_256), .ZN(n_1_241));
   INV_X1 i_1_426 (.A(n_1_242), .ZN(n_167));
   AOI222_X1 i_1_427 (.A1(\temp2[2] [20]), .A2(n_1_257), .B1(\temp1[2] [20]), 
      .B2(n_1_258), .C1(n_183), .C2(n_1_256), .ZN(n_1_242));
   INV_X1 i_1_428 (.A(n_1_243), .ZN(n_168));
   AOI222_X1 i_1_429 (.A1(\temp2[2] [21]), .A2(n_1_257), .B1(\temp1[2] [21]), 
      .B2(n_1_258), .C1(n_184), .C2(n_1_256), .ZN(n_1_243));
   INV_X1 i_1_430 (.A(n_1_244), .ZN(n_169));
   AOI222_X1 i_1_431 (.A1(\temp2[2] [22]), .A2(n_1_257), .B1(\temp1[2] [22]), 
      .B2(n_1_258), .C1(n_185), .C2(n_1_256), .ZN(n_1_244));
   INV_X1 i_1_432 (.A(n_1_245), .ZN(n_170));
   AOI222_X1 i_1_433 (.A1(\temp2[2] [23]), .A2(n_1_257), .B1(\temp1[2] [23]), 
      .B2(n_1_258), .C1(n_186), .C2(n_1_256), .ZN(n_1_245));
   INV_X1 i_1_434 (.A(n_1_246), .ZN(n_171));
   AOI222_X1 i_1_435 (.A1(\temp2[2] [24]), .A2(n_1_257), .B1(\temp1[2] [24]), 
      .B2(n_1_258), .C1(n_187), .C2(n_1_256), .ZN(n_1_246));
   INV_X1 i_1_436 (.A(n_1_247), .ZN(n_172));
   AOI222_X1 i_1_437 (.A1(\temp2[2] [25]), .A2(n_1_257), .B1(\temp1[2] [25]), 
      .B2(n_1_258), .C1(n_188), .C2(n_1_256), .ZN(n_1_247));
   INV_X1 i_1_438 (.A(n_1_248), .ZN(n_173));
   AOI222_X1 i_1_439 (.A1(\temp2[2] [26]), .A2(n_1_257), .B1(\temp1[2] [26]), 
      .B2(n_1_258), .C1(n_189), .C2(n_1_256), .ZN(n_1_248));
   INV_X1 i_1_440 (.A(n_1_249), .ZN(n_174));
   AOI222_X1 i_1_441 (.A1(\temp2[2] [27]), .A2(n_1_257), .B1(\temp1[2] [27]), 
      .B2(n_1_258), .C1(n_190), .C2(n_1_256), .ZN(n_1_249));
   INV_X1 i_1_442 (.A(n_1_250), .ZN(n_175));
   AOI222_X1 i_1_443 (.A1(\temp2[2] [28]), .A2(n_1_257), .B1(\temp1[2] [28]), 
      .B2(n_1_258), .C1(n_191), .C2(n_1_256), .ZN(n_1_250));
   INV_X1 i_1_444 (.A(n_1_251), .ZN(n_176));
   AOI222_X1 i_1_445 (.A1(\temp2[2] [29]), .A2(n_1_257), .B1(\temp1[2] [29]), 
      .B2(n_1_258), .C1(n_192), .C2(n_1_256), .ZN(n_1_251));
   INV_X1 i_1_446 (.A(n_1_252), .ZN(n_177));
   AOI222_X1 i_1_447 (.A1(\temp2[2] [30]), .A2(n_1_257), .B1(\temp1[2] [30]), 
      .B2(n_1_258), .C1(n_193), .C2(n_1_256), .ZN(n_1_252));
   INV_X1 i_1_448 (.A(n_1_253), .ZN(n_178));
   AOI221_X1 i_1_449 (.A(n_1_255), .B1(\temp1[2] [31]), .B2(n_1_258), .C1(
      \temp2[2] [31]), .C2(n_1_257), .ZN(n_1_253));
   INV_X1 i_1_450 (.A(n_1_254), .ZN(n_179));
   AOI221_X1 i_1_451 (.A(n_1_255), .B1(\temp1[2] [32]), .B2(n_1_258), .C1(
      \temp2[2] [32]), .C2(n_1_257), .ZN(n_1_254));
   AND2_X1 i_1_452 (.A1(n_194), .A2(n_1_256), .ZN(n_1_255));
   NOR2_X1 i_1_453 (.A1(n_1_258), .A2(n_1_257), .ZN(n_1_256));
   NOR2_X1 i_1_454 (.A1(n_1_16), .A2(r[1]), .ZN(n_1_257));
   NOR2_X1 i_1_455 (.A1(r[2]), .A2(n_1_15), .ZN(n_1_258));
   INV_X1 i_1_456 (.A(n_1_259), .ZN(n_180));
   AOI222_X1 i_1_457 (.A1(\temp1[1] [18]), .A2(n_1_13), .B1(r[1]), .B2(n_196), 
      .C1(\temp2[1] [18]), .C2(n_1_274), .ZN(n_1_259));
   INV_X1 i_1_458 (.A(n_1_260), .ZN(n_181));
   AOI222_X1 i_1_459 (.A1(mn[3]), .A2(n_1_12), .B1(\temp2[1] [19]), .B2(n_1_274), 
      .C1(\temp1[1] [19]), .C2(n_1_13), .ZN(n_1_260));
   INV_X1 i_1_460 (.A(n_1_261), .ZN(n_182));
   AOI222_X1 i_1_461 (.A1(mn[4]), .A2(n_1_12), .B1(\temp2[1] [20]), .B2(n_1_274), 
      .C1(\temp1[1] [20]), .C2(n_1_13), .ZN(n_1_261));
   INV_X1 i_1_462 (.A(n_1_262), .ZN(n_183));
   AOI222_X1 i_1_463 (.A1(mn[5]), .A2(n_1_12), .B1(\temp2[1] [21]), .B2(n_1_274), 
      .C1(\temp1[1] [21]), .C2(n_1_13), .ZN(n_1_262));
   INV_X1 i_1_464 (.A(n_1_263), .ZN(n_184));
   AOI222_X1 i_1_465 (.A1(mn[6]), .A2(n_1_12), .B1(\temp2[1] [22]), .B2(n_1_274), 
      .C1(\temp1[1] [22]), .C2(n_1_13), .ZN(n_1_263));
   INV_X1 i_1_466 (.A(n_1_264), .ZN(n_185));
   AOI222_X1 i_1_467 (.A1(mn[7]), .A2(n_1_12), .B1(\temp2[1] [23]), .B2(n_1_274), 
      .C1(\temp1[1] [23]), .C2(n_1_13), .ZN(n_1_264));
   INV_X1 i_1_468 (.A(n_1_265), .ZN(n_186));
   AOI222_X1 i_1_469 (.A1(mn[8]), .A2(n_1_12), .B1(\temp2[1] [24]), .B2(n_1_274), 
      .C1(\temp1[1] [24]), .C2(n_1_13), .ZN(n_1_265));
   INV_X1 i_1_470 (.A(n_1_266), .ZN(n_187));
   AOI222_X1 i_1_471 (.A1(mn[9]), .A2(n_1_12), .B1(\temp2[1] [25]), .B2(n_1_274), 
      .C1(\temp1[1] [25]), .C2(n_1_13), .ZN(n_1_266));
   INV_X1 i_1_472 (.A(n_1_267), .ZN(n_188));
   AOI222_X1 i_1_473 (.A1(mn[10]), .A2(n_1_12), .B1(\temp2[1] [26]), .B2(n_1_274), 
      .C1(\temp1[1] [26]), .C2(n_1_13), .ZN(n_1_267));
   INV_X1 i_1_474 (.A(n_1_268), .ZN(n_189));
   AOI222_X1 i_1_475 (.A1(r[1]), .A2(n_205), .B1(\temp2[1] [27]), .B2(n_1_274), 
      .C1(\temp1[1] [27]), .C2(n_1_13), .ZN(n_1_268));
   INV_X1 i_1_476 (.A(n_1_269), .ZN(n_190));
   AOI222_X1 i_1_477 (.A1(r[1]), .A2(n_206), .B1(\temp2[1] [28]), .B2(n_1_274), 
      .C1(\temp1[1] [28]), .C2(n_1_13), .ZN(n_1_269));
   INV_X1 i_1_478 (.A(n_1_270), .ZN(n_191));
   AOI222_X1 i_1_479 (.A1(r[1]), .A2(n_207), .B1(\temp2[1] [29]), .B2(n_1_274), 
      .C1(\temp1[1] [29]), .C2(n_1_13), .ZN(n_1_270));
   INV_X1 i_1_480 (.A(n_1_271), .ZN(n_192));
   AOI222_X1 i_1_481 (.A1(r[1]), .A2(n_208), .B1(\temp2[1] [30]), .B2(n_1_274), 
      .C1(\temp1[1] [30]), .C2(n_1_13), .ZN(n_1_271));
   INV_X1 i_1_482 (.A(n_1_272), .ZN(n_193));
   AOI221_X1 i_1_483 (.A(n_1_275), .B1(\temp2[1] [31]), .B2(n_1_274), .C1(
      \temp1[1] [31]), .C2(n_1_13), .ZN(n_1_272));
   INV_X1 i_1_484 (.A(n_1_273), .ZN(n_194));
   AOI221_X1 i_1_485 (.A(n_1_275), .B1(\temp2[1] [32]), .B2(n_1_274), .C1(
      \temp1[1] [32]), .C2(n_1_13), .ZN(n_1_273));
   NOR2_X1 i_1_486 (.A1(n_1_15), .A2(r[0]), .ZN(n_1_274));
   AND2_X1 i_1_487 (.A1(mn[15]), .A2(n_1_12), .ZN(n_1_275));
   NOR2_X1 i_1_488 (.A1(n_1_15), .A2(n_1_14), .ZN(n_1_12));
   NOR2_X1 i_1_489 (.A1(r[1]), .A2(n_1_14), .ZN(n_1_13));
   AND2_X1 i_1_490 (.A1(r[0]), .A2(mn[1]), .ZN(n_195));
   AND2_X1 i_1_491 (.A1(r[0]), .A2(mn[2]), .ZN(n_196));
   AND2_X1 i_1_492 (.A1(r[0]), .A2(mn[3]), .ZN(n_197));
   AND2_X1 i_1_493 (.A1(r[0]), .A2(mn[4]), .ZN(n_198));
   AND2_X1 i_1_494 (.A1(r[0]), .A2(mn[5]), .ZN(n_199));
   AND2_X1 i_1_495 (.A1(r[0]), .A2(mn[6]), .ZN(n_200));
   AND2_X1 i_1_496 (.A1(r[0]), .A2(mn[7]), .ZN(n_201));
   AND2_X1 i_1_497 (.A1(r[0]), .A2(mn[8]), .ZN(n_202));
   AND2_X1 i_1_498 (.A1(r[0]), .A2(mn[9]), .ZN(n_203));
   AND2_X1 i_1_499 (.A1(r[0]), .A2(mn[10]), .ZN(n_204));
   AND2_X1 i_1_500 (.A1(r[0]), .A2(mn[11]), .ZN(n_205));
   AND2_X1 i_1_501 (.A1(r[0]), .A2(mn[12]), .ZN(n_206));
   AND2_X1 i_1_502 (.A1(r[0]), .A2(mn[13]), .ZN(n_207));
   AND2_X1 i_1_503 (.A1(r[0]), .A2(mn[14]), .ZN(n_208));
   AND2_X1 i_1_504 (.A1(r[0]), .A2(mn[15]), .ZN(n_209));
   INV_X1 i_1_505 (.A(r[0]), .ZN(n_1_14));
   INV_X1 i_1_506 (.A(r[1]), .ZN(n_1_15));
   INV_X1 i_1_507 (.A(r[2]), .ZN(n_1_16));
   INV_X1 i_1_508 (.A(r[3]), .ZN(n_1_17));
   INV_X1 i_1_509 (.A(r[4]), .ZN(n_1_18));
   INV_X1 i_1_510 (.A(r[5]), .ZN(n_1_19));
   INV_X1 i_1_511 (.A(r[6]), .ZN(n_1_20));
   INV_X1 i_1_512 (.A(r[7]), .ZN(n_1_21));
   INV_X1 i_1_513 (.A(r[8]), .ZN(n_1_22));
   INV_X1 i_1_514 (.A(r[9]), .ZN(n_1_23));
   INV_X1 i_1_515 (.A(r[10]), .ZN(n_1_24));
   INV_X1 i_1_516 (.A(r[11]), .ZN(n_1_25));
   INV_X1 i_1_517 (.A(r[12]), .ZN(n_1_26));
   INV_X1 i_1_518 (.A(r[13]), .ZN(n_1_27));
endmodule

module reg__3_24(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;

   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_13), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_13), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_13), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_13), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_13), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_13), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_13), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_13), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_13), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_13), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_13), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_13), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_13), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_14), .B1(n_0_13), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_14), .B1(n_0_13), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_14), .B1(n_0_13), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_14), .B1(n_0_13), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_14), .B1(n_0_13), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_14), .B1(n_0_13), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_14), .B1(n_0_13), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_14), .B1(n_0_13), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_14), .B1(n_0_13), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_14), .B1(n_0_13), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_14), .B1(n_0_13), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_14), .B1(n_0_13), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_14), .B1(n_0_13), .B2(Q[12]), .ZN(n_0_12));
   NOR2_X1 i_0_26 (.A1(rst), .A2(load), .ZN(n_0_13));
   NOR2_X1 i_0_27 (.A1(n_0_15), .A2(rst), .ZN(n_0_14));
   INV_X1 i_0_28 (.A(load), .ZN(n_0_15));
   INV_X1 i_0_29 (.A(Clk), .ZN(n_13));
endmodule

module Decoder1(s, firstRaw, d);
   input [2:0]s;
   input firstRaw;
   output [1:10]d;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   AND3_X1 i_0_0 (.A1(s[2]), .A2(s[1]), .A3(s[0]), .ZN(d[10]));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(d[9]));
   AOI21_X1 i_0_2 (.A(d[1]), .B1(s[1]), .B2(s[2]), .ZN(n_0_0));
   AND2_X1 i_0_3 (.A1(firstRaw), .A2(d[4]), .ZN(d[8]));
   NOR3_X1 i_0_4 (.A1(n_0_1), .A2(s[0]), .A3(firstRaw), .ZN(d[7]));
   NOR3_X1 i_0_5 (.A1(n_0_3), .A2(n_0_2), .A3(s[2]), .ZN(d[6]));
   AOI21_X1 i_0_6 (.A(n_0_1), .B1(n_0_2), .B2(firstRaw), .ZN(d[5]));
   NOR2_X1 i_0_7 (.A1(n_0_1), .A2(s[0]), .ZN(d[4]));
   NAND2_X1 i_0_8 (.A1(n_0_3), .A2(s[2]), .ZN(n_0_1));
   NOR3_X1 i_0_9 (.A1(n_0_2), .A2(s[1]), .A3(s[2]), .ZN(d[1]));
   INV_X1 i_0_10 (.A(s[0]), .ZN(n_0_2));
   INV_X1 i_0_11 (.A(s[1]), .ZN(n_0_3));
endmodule

module reg__3_44(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module twoInpMux(In0, In1, selector, out1);
   input [15:0]In0;
   input [15:0]In1;
   input selector;
   output [15:0]out1;

   MUX2_X1 i_0_0 (.A(In0[0]), .B(In1[0]), .S(selector), .Z(out1[0]));
   MUX2_X1 i_0_1 (.A(In0[1]), .B(In1[1]), .S(selector), .Z(out1[1]));
   MUX2_X1 i_0_2 (.A(In0[2]), .B(In1[2]), .S(selector), .Z(out1[2]));
   MUX2_X1 i_0_3 (.A(In0[3]), .B(In1[3]), .S(selector), .Z(out1[3]));
   MUX2_X1 i_0_4 (.A(In0[4]), .B(In1[4]), .S(selector), .Z(out1[4]));
   MUX2_X1 i_0_5 (.A(In0[5]), .B(In1[5]), .S(selector), .Z(out1[5]));
   MUX2_X1 i_0_6 (.A(In0[6]), .B(In1[6]), .S(selector), .Z(out1[6]));
   MUX2_X1 i_0_7 (.A(In0[7]), .B(In1[7]), .S(selector), .Z(out1[7]));
   MUX2_X1 i_0_8 (.A(In0[8]), .B(In1[8]), .S(selector), .Z(out1[8]));
   MUX2_X1 i_0_9 (.A(In0[9]), .B(In1[9]), .S(selector), .Z(out1[9]));
   MUX2_X1 i_0_10 (.A(In0[10]), .B(In1[10]), .S(selector), .Z(out1[10]));
   MUX2_X1 i_0_11 (.A(In0[11]), .B(In1[11]), .S(selector), .Z(out1[11]));
   MUX2_X1 i_0_12 (.A(In0[12]), .B(In1[12]), .S(selector), .Z(out1[12]));
   MUX2_X1 i_0_13 (.A(In0[13]), .B(In1[13]), .S(selector), .Z(out1[13]));
   MUX2_X1 i_0_14 (.A(In0[14]), .B(In1[14]), .S(selector), .Z(out1[14]));
   MUX2_X1 i_0_15 (.A(In0[15]), .B(In1[15]), .S(selector), .Z(out1[15]));
endmodule

module reg__3_64(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module M1Add1Mux(Init, E, Ti, A, Xstore, XS1, XS2, selector, Var1, Var2, Var3, 
      Add);
   input [15:0]Init;
   input [15:0]E;
   input [15:0]Ti;
   input [15:0]A;
   input [15:0]Xstore;
   input [15:0]XS1;
   input [15:0]XS2;
   input [2:0]selector;
   input Var1;
   input Var2;
   input Var3;
   output [15:0]Add;

   wire n_0_0;
   wire n_0_2;
   wire n_0_4;
   wire n_0_6;
   wire n_0_8;
   wire n_0_10;
   wire n_0_12;
   wire n_0_14;
   wire n_0_16;
   wire n_0_18;
   wire n_0_20;
   wire n_0_22;
   wire n_0_24;
   wire n_0_26;
   wire n_0_28;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_35;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_1;
   wire n_0_34;
   wire n_0_29;
   wire n_0_27;
   wire n_0_25;
   wire n_0_23;
   wire n_0_21;
   wire n_0_19;
   wire n_0_17;
   wire n_0_15;
   wire n_0_13;
   wire n_0_11;
   wire n_0_9;
   wire n_0_7;
   wire n_0_5;
   wire n_0_3;
   wire n_0_36;

   NAND2_X1 i_0_0 (.A1(n_0_36), .A2(n_0_0), .ZN(Add[0]));
   AOI22_X1 i_0_1 (.A1(Xstore[0]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[0]), 
      .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_2), .ZN(Add[1]));
   AOI22_X1 i_0_4 (.A1(Xstore[1]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[1]), 
      .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(n_0_5), .A2(n_0_4), .ZN(Add[2]));
   AOI22_X1 i_0_7 (.A1(Xstore[2]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[2]), 
      .ZN(n_0_4));
   NAND2_X1 i_0_9 (.A1(n_0_7), .A2(n_0_6), .ZN(Add[3]));
   AOI22_X1 i_0_10 (.A1(Xstore[3]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[3]), 
      .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(n_0_9), .A2(n_0_8), .ZN(Add[4]));
   AOI22_X1 i_0_13 (.A1(Xstore[4]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[4]), 
      .ZN(n_0_8));
   NAND2_X1 i_0_15 (.A1(n_0_11), .A2(n_0_10), .ZN(Add[5]));
   AOI22_X1 i_0_16 (.A1(Xstore[5]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[5]), 
      .ZN(n_0_10));
   NAND2_X1 i_0_18 (.A1(n_0_13), .A2(n_0_12), .ZN(Add[6]));
   AOI22_X1 i_0_19 (.A1(Xstore[6]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[6]), 
      .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(n_0_15), .A2(n_0_14), .ZN(Add[7]));
   AOI22_X1 i_0_22 (.A1(Xstore[7]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[7]), 
      .ZN(n_0_14));
   NAND2_X1 i_0_24 (.A1(n_0_17), .A2(n_0_16), .ZN(Add[8]));
   AOI22_X1 i_0_25 (.A1(Xstore[8]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[8]), 
      .ZN(n_0_16));
   NAND2_X1 i_0_27 (.A1(n_0_19), .A2(n_0_18), .ZN(Add[9]));
   AOI22_X1 i_0_28 (.A1(Xstore[9]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[9]), 
      .ZN(n_0_18));
   NAND2_X1 i_0_30 (.A1(n_0_21), .A2(n_0_20), .ZN(Add[10]));
   AOI22_X1 i_0_31 (.A1(Xstore[10]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[10]), 
      .ZN(n_0_20));
   NAND2_X1 i_0_33 (.A1(n_0_23), .A2(n_0_22), .ZN(Add[11]));
   AOI22_X1 i_0_34 (.A1(Xstore[11]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[11]), 
      .ZN(n_0_22));
   NAND2_X1 i_0_36 (.A1(n_0_25), .A2(n_0_24), .ZN(Add[12]));
   AOI22_X1 i_0_37 (.A1(Xstore[12]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[12]), 
      .ZN(n_0_24));
   NAND2_X1 i_0_39 (.A1(n_0_27), .A2(n_0_26), .ZN(Add[13]));
   AOI22_X1 i_0_40 (.A1(Xstore[13]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[13]), 
      .ZN(n_0_26));
   NAND2_X1 i_0_42 (.A1(n_0_29), .A2(n_0_28), .ZN(Add[14]));
   AOI22_X1 i_0_43 (.A1(Xstore[14]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[14]), 
      .ZN(n_0_28));
   NAND2_X1 i_0_45 (.A1(n_0_34), .A2(n_0_30), .ZN(Add[15]));
   AOI22_X1 i_0_46 (.A1(Xstore[15]), .A2(n_0_32), .B1(n_0_31), .B2(XS2[15]), 
      .ZN(n_0_30));
   NOR2_X1 i_0_47 (.A1(n_0_1), .A2(n_0_33), .ZN(n_0_31));
   NOR2_X1 i_0_48 (.A1(n_0_33), .A2(Var2), .ZN(n_0_32));
   OR4_X1 i_0_49 (.A1(n_0_40), .A2(selector[0]), .A3(Var1), .A4(Var3), .ZN(
      n_0_33));
   NOR3_X1 i_0_50 (.A1(n_0_41), .A2(selector[1]), .A3(selector[0]), .ZN(n_0_35));
   NOR2_X1 i_0_51 (.A1(n_0_38), .A2(n_0_40), .ZN(n_0_37));
   AOI21_X1 i_0_52 (.A(selector[0]), .B1(n_0_39), .B2(Var1), .ZN(n_0_38));
   NOR2_X1 i_0_53 (.A1(Var3), .A2(Var2), .ZN(n_0_39));
   NAND2_X1 i_0_54 (.A1(selector[2]), .A2(selector[1]), .ZN(n_0_40));
   INV_X1 i_0_55 (.A(selector[2]), .ZN(n_0_41));
   INV_X1 i_0_56 (.A(Var2), .ZN(n_0_1));
   AOI22_X1 i_0_2 (.A1(XS1[15]), .A2(n_0_37), .B1(n_0_35), .B2(A[15]), .ZN(
      n_0_34));
   AOI22_X1 i_0_5 (.A1(XS1[14]), .A2(n_0_37), .B1(n_0_35), .B2(A[14]), .ZN(
      n_0_29));
   AOI22_X1 i_0_8 (.A1(XS1[13]), .A2(n_0_37), .B1(n_0_35), .B2(A[13]), .ZN(
      n_0_27));
   AOI22_X1 i_0_11 (.A1(XS1[12]), .A2(n_0_37), .B1(n_0_35), .B2(A[12]), .ZN(
      n_0_25));
   AOI22_X1 i_0_14 (.A1(XS1[11]), .A2(n_0_37), .B1(n_0_35), .B2(A[11]), .ZN(
      n_0_23));
   AOI22_X1 i_0_17 (.A1(XS1[10]), .A2(n_0_37), .B1(n_0_35), .B2(A[10]), .ZN(
      n_0_21));
   AOI22_X1 i_0_20 (.A1(XS1[9]), .A2(n_0_37), .B1(n_0_35), .B2(A[9]), .ZN(n_0_19));
   AOI22_X1 i_0_23 (.A1(XS1[8]), .A2(n_0_37), .B1(n_0_35), .B2(A[8]), .ZN(n_0_17));
   AOI22_X1 i_0_26 (.A1(XS1[7]), .A2(n_0_37), .B1(n_0_35), .B2(A[7]), .ZN(n_0_15));
   AOI22_X1 i_0_29 (.A1(XS1[6]), .A2(n_0_37), .B1(n_0_35), .B2(A[6]), .ZN(n_0_13));
   AOI22_X1 i_0_32 (.A1(XS1[5]), .A2(n_0_37), .B1(n_0_35), .B2(A[5]), .ZN(n_0_11));
   AOI22_X1 i_0_35 (.A1(XS1[4]), .A2(n_0_37), .B1(n_0_35), .B2(A[4]), .ZN(n_0_9));
   AOI22_X1 i_0_38 (.A1(XS1[3]), .A2(n_0_37), .B1(n_0_35), .B2(A[3]), .ZN(n_0_7));
   AOI22_X1 i_0_41 (.A1(XS1[2]), .A2(n_0_37), .B1(n_0_35), .B2(A[2]), .ZN(n_0_5));
   AOI22_X1 i_0_44 (.A1(XS1[1]), .A2(n_0_37), .B1(n_0_35), .B2(A[1]), .ZN(n_0_3));
   AOI22_X1 i_0_57 (.A1(XS1[0]), .A2(n_0_37), .B1(n_0_35), .B2(A[0]), .ZN(n_0_36));
endmodule

module M1Add2Mux(H, Xn, Xprev, Xs2, selector, Add);
   input [15:0]H;
   input [15:0]Xn;
   input [15:0]Xprev;
   input [15:0]Xs2;
   input [2:0]selector;
   output [15:0]Add;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;

   OAI21_X1 i_0_0 (.A(n_0_0), .B1(n_0_1), .B2(selector[0]), .ZN(Add[0]));
   AOI22_X1 i_0_1 (.A1(Xn[0]), .A2(n_0_19), .B1(n_0_18), .B2(Xs2[0]), .ZN(n_0_0));
   OAI21_X1 i_0_2 (.A(selector[1]), .B1(n_0_21), .B2(Xprev[0]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(Add[1]));
   AOI222_X1 i_0_4 (.A1(Xs2[1]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[1]), 
      .C1(Xn[1]), .C2(n_0_19), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_3), .ZN(Add[2]));
   AOI222_X1 i_0_6 (.A1(Xs2[2]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[2]), 
      .C1(Xn[2]), .C2(n_0_19), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_4), .ZN(Add[3]));
   AOI222_X1 i_0_8 (.A1(Xs2[3]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[3]), 
      .C1(Xn[3]), .C2(n_0_19), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(Add[4]));
   AOI222_X1 i_0_10 (.A1(Xs2[4]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[4]), 
      .C1(Xn[4]), .C2(n_0_19), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_6), .ZN(Add[5]));
   AOI222_X1 i_0_12 (.A1(Xs2[5]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[5]), 
      .C1(Xn[5]), .C2(n_0_19), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_7), .ZN(Add[6]));
   AOI222_X1 i_0_14 (.A1(Xs2[6]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[6]), 
      .C1(Xn[6]), .C2(n_0_19), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_8), .ZN(Add[7]));
   AOI222_X1 i_0_16 (.A1(Xs2[7]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[7]), 
      .C1(Xn[7]), .C2(n_0_19), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_9), .ZN(Add[8]));
   AOI222_X1 i_0_18 (.A1(Xs2[8]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[8]), 
      .C1(Xn[8]), .C2(n_0_19), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_10), .ZN(Add[9]));
   AOI222_X1 i_0_20 (.A1(Xs2[9]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[9]), 
      .C1(Xn[9]), .C2(n_0_19), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_11), .ZN(Add[10]));
   AOI222_X1 i_0_22 (.A1(Xs2[10]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[10]), 
      .C1(Xn[10]), .C2(n_0_19), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_12), .ZN(Add[11]));
   AOI222_X1 i_0_24 (.A1(Xs2[11]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[11]), 
      .C1(Xn[11]), .C2(n_0_19), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_13), .ZN(Add[12]));
   AOI222_X1 i_0_26 (.A1(Xs2[12]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[12]), 
      .C1(Xn[12]), .C2(n_0_19), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_14), .ZN(Add[13]));
   AOI222_X1 i_0_28 (.A1(Xs2[13]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[13]), 
      .C1(Xn[13]), .C2(n_0_19), .ZN(n_0_14));
   INV_X1 i_0_29 (.A(n_0_15), .ZN(Add[14]));
   AOI222_X1 i_0_30 (.A1(Xs2[14]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[14]), 
      .C1(Xn[14]), .C2(n_0_19), .ZN(n_0_15));
   INV_X1 i_0_31 (.A(n_0_16), .ZN(Add[15]));
   AOI222_X1 i_0_32 (.A1(Xs2[15]), .A2(n_0_18), .B1(n_0_17), .B2(Xprev[15]), 
      .C1(Xn[15]), .C2(n_0_19), .ZN(n_0_16));
   NOR3_X1 i_0_33 (.A1(n_0_21), .A2(n_0_20), .A3(selector[0]), .ZN(n_0_17));
   AND3_X1 i_0_34 (.A1(selector[2]), .A2(selector[1]), .A3(selector[0]), 
      .ZN(n_0_18));
   NOR3_X1 i_0_35 (.A1(n_0_21), .A2(selector[1]), .A3(selector[0]), .ZN(n_0_19));
   INV_X1 i_0_36 (.A(selector[1]), .ZN(n_0_20));
   INV_X1 i_0_37 (.A(selector[2]), .ZN(n_0_21));
endmodule

module M2Add1Mux(Ucalc, Un, Ustore, selector, firstRaw, Add);
   input [15:0]Ucalc;
   input [15:0]Un;
   input [15:0]Ustore;
   input [2:0]selector;
   input firstRaw;
   output [15:0]Add;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(Add[0]));
   AOI22_X1 i_0_1 (.A1(Un[0]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[0]), .ZN(
      n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(Add[1]));
   AOI22_X1 i_0_3 (.A1(Un[1]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[1]), .ZN(
      n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(Add[2]));
   AOI22_X1 i_0_5 (.A1(Un[2]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[2]), .ZN(
      n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(Add[3]));
   AOI22_X1 i_0_7 (.A1(Un[3]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[3]), .ZN(
      n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(Add[4]));
   AOI22_X1 i_0_9 (.A1(Un[4]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[4]), .ZN(
      n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(Add[5]));
   AOI22_X1 i_0_11 (.A1(Un[5]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[5]), 
      .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(Add[6]));
   AOI22_X1 i_0_13 (.A1(Un[6]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[6]), 
      .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(Add[7]));
   AOI22_X1 i_0_15 (.A1(Un[7]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[7]), 
      .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(Add[8]));
   AOI22_X1 i_0_17 (.A1(Un[8]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[8]), 
      .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(Add[9]));
   AOI22_X1 i_0_19 (.A1(Un[9]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[9]), 
      .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(Add[10]));
   AOI22_X1 i_0_21 (.A1(Un[10]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[10]), 
      .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(Add[11]));
   AOI22_X1 i_0_23 (.A1(Un[11]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[11]), 
      .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(Add[12]));
   AOI22_X1 i_0_25 (.A1(Un[12]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[12]), 
      .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(Add[13]));
   AOI22_X1 i_0_27 (.A1(Un[13]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[13]), 
      .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(Add[14]));
   AOI22_X1 i_0_29 (.A1(Un[14]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[14]), 
      .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(Add[15]));
   AOI22_X1 i_0_31 (.A1(Un[15]), .A2(n_0_17), .B1(n_0_16), .B2(Ucalc[15]), 
      .ZN(n_0_15));
   NOR3_X1 i_0_32 (.A1(n_0_18), .A2(n_0_19), .A3(selector[1]), .ZN(n_0_16));
   NOR4_X1 i_0_33 (.A1(n_0_20), .A2(n_0_19), .A3(selector[1]), .A4(selector[0]), 
      .ZN(n_0_17));
   NOR2_X1 i_0_34 (.A1(n_0_20), .A2(selector[0]), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(selector[2]), .ZN(n_0_19));
   INV_X1 i_0_36 (.A(firstRaw), .ZN(n_0_20));
endmodule

module M2Add2Mux(B, Uz, selector, firstRaw, Add);
   input [15:0]B;
   input [15:0]Uz;
   input [2:0]selector;
   input firstRaw;
   output [15:0]Add;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   INV_X1 i_0_0 (.A(selector[2]), .ZN(n_0_0));
   NOR4_X1 i_0_1 (.A1(n_0_0), .A2(firstRaw), .A3(selector[0]), .A4(selector[1]), 
      .ZN(n_0_1));
   NOR4_X1 i_0_2 (.A1(n_0_1), .A2(n_0_0), .A3(selector[0]), .A4(selector[1]), 
      .ZN(n_0_2));
   AOI22_X1 i_0_3 (.A1(n_0_2), .A2(Uz[0]), .B1(n_0_1), .B2(B[0]), .ZN(n_0_3));
   INV_X1 i_0_4 (.A(n_0_3), .ZN(Add[0]));
   AOI22_X1 i_0_5 (.A1(n_0_2), .A2(Uz[1]), .B1(n_0_1), .B2(B[1]), .ZN(n_0_4));
   INV_X1 i_0_6 (.A(n_0_4), .ZN(Add[1]));
   AOI22_X1 i_0_7 (.A1(n_0_2), .A2(Uz[2]), .B1(n_0_1), .B2(B[2]), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(n_0_5), .ZN(Add[2]));
   AOI22_X1 i_0_9 (.A1(n_0_2), .A2(Uz[3]), .B1(n_0_1), .B2(B[3]), .ZN(n_0_6));
   INV_X1 i_0_10 (.A(n_0_6), .ZN(Add[3]));
   AOI22_X1 i_0_11 (.A1(n_0_2), .A2(Uz[4]), .B1(n_0_1), .B2(B[4]), .ZN(n_0_7));
   INV_X1 i_0_12 (.A(n_0_7), .ZN(Add[4]));
   AOI22_X1 i_0_13 (.A1(n_0_2), .A2(Uz[5]), .B1(n_0_1), .B2(B[5]), .ZN(n_0_8));
   INV_X1 i_0_14 (.A(n_0_8), .ZN(Add[5]));
   AOI22_X1 i_0_15 (.A1(n_0_2), .A2(Uz[6]), .B1(n_0_1), .B2(B[6]), .ZN(n_0_9));
   INV_X1 i_0_16 (.A(n_0_9), .ZN(Add[6]));
   AOI22_X1 i_0_17 (.A1(n_0_2), .A2(Uz[7]), .B1(n_0_1), .B2(B[7]), .ZN(n_0_10));
   INV_X1 i_0_18 (.A(n_0_10), .ZN(Add[7]));
   AOI22_X1 i_0_19 (.A1(n_0_2), .A2(Uz[8]), .B1(n_0_1), .B2(B[8]), .ZN(n_0_11));
   INV_X1 i_0_20 (.A(n_0_11), .ZN(Add[8]));
   AOI22_X1 i_0_21 (.A1(n_0_2), .A2(Uz[9]), .B1(n_0_1), .B2(B[9]), .ZN(n_0_12));
   INV_X1 i_0_22 (.A(n_0_12), .ZN(Add[9]));
   AOI22_X1 i_0_23 (.A1(n_0_2), .A2(Uz[10]), .B1(n_0_1), .B2(B[10]), .ZN(n_0_13));
   INV_X1 i_0_24 (.A(n_0_13), .ZN(Add[10]));
   AOI22_X1 i_0_25 (.A1(n_0_2), .A2(Uz[11]), .B1(n_0_1), .B2(B[11]), .ZN(n_0_14));
   INV_X1 i_0_26 (.A(n_0_14), .ZN(Add[11]));
   AOI22_X1 i_0_27 (.A1(n_0_2), .A2(Uz[12]), .B1(n_0_1), .B2(B[12]), .ZN(n_0_15));
   INV_X1 i_0_28 (.A(n_0_15), .ZN(Add[12]));
   AOI22_X1 i_0_29 (.A1(n_0_2), .A2(Uz[13]), .B1(n_0_1), .B2(B[13]), .ZN(n_0_16));
   INV_X1 i_0_30 (.A(n_0_16), .ZN(Add[13]));
   AOI22_X1 i_0_31 (.A1(n_0_2), .A2(Uz[14]), .B1(n_0_1), .B2(B[14]), .ZN(n_0_17));
   INV_X1 i_0_32 (.A(n_0_17), .ZN(Add[14]));
   AOI22_X1 i_0_33 (.A1(n_0_2), .A2(Uz[15]), .B1(n_0_1), .B2(B[15]), .ZN(n_0_18));
   INV_X1 i_0_34 (.A(n_0_18), .ZN(Add[15]));
endmodule

module reg__3_84(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module reg__3_104(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;

   DFF_X1 \Q_reg[15]  (.D(n_15), .CK(n_16), .Q(Q[15]), .QN());
   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_16), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_16), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_16), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_16), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_16), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_16), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_16), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_16), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_16), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_16), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_16), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_16), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_16), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_16), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_16), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_17), .B1(n_0_16), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_17), .B1(n_0_16), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_17), .B1(n_0_16), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_17), .B1(n_0_16), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_17), .B1(n_0_16), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_17), .B1(n_0_16), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_17), .B1(n_0_16), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_17), .B1(n_0_16), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_17), .B1(n_0_16), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_17), .B1(n_0_16), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_17), .B1(n_0_16), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_17), .B1(n_0_16), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_17), .B1(n_0_16), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_17), .B1(n_0_16), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_17), .B1(n_0_16), .B2(Q[14]), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_15));
   AOI22_X1 i_0_31 (.A1(D[15]), .A2(n_0_17), .B1(n_0_16), .B2(Q[15]), .ZN(n_0_15));
   NOR2_X1 i_0_32 (.A1(rst), .A2(load), .ZN(n_0_16));
   NOR2_X1 i_0_33 (.A1(n_0_18), .A2(rst), .ZN(n_0_17));
   INV_X1 i_0_34 (.A(load), .ZN(n_0_18));
   INV_X1 i_0_35 (.A(Clk), .ZN(n_16));
endmodule

module reg__3_124(D, load, Clk, Q, rst);
   input [15:0]D;
   input load;
   input Clk;
   output [15:0]Q;
   input rst;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;

   DFF_X1 \Q_reg[14]  (.D(n_14), .CK(n_15), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[13]  (.D(n_13), .CK(n_15), .Q(Q[13]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_12), .CK(n_15), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_11), .CK(n_15), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_10), .CK(n_15), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_9), .CK(n_15), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_8), .CK(n_15), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_7), .CK(n_15), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_6), .CK(n_15), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_5), .CK(n_15), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_4), .CK(n_15), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_3), .CK(n_15), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_2), .CK(n_15), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_1), .CK(n_15), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0), .CK(n_15), .Q(Q[0]), .QN());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(n_0));
   AOI22_X1 i_0_1 (.A1(D[0]), .A2(n_0_16), .B1(n_0_15), .B2(Q[0]), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_1));
   AOI22_X1 i_0_3 (.A1(D[1]), .A2(n_0_16), .B1(n_0_15), .B2(Q[1]), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_2));
   AOI22_X1 i_0_5 (.A1(D[2]), .A2(n_0_16), .B1(n_0_15), .B2(Q[2]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_3));
   AOI22_X1 i_0_7 (.A1(D[3]), .A2(n_0_16), .B1(n_0_15), .B2(Q[3]), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_4));
   AOI22_X1 i_0_9 (.A1(D[4]), .A2(n_0_16), .B1(n_0_15), .B2(Q[4]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_5));
   AOI22_X1 i_0_11 (.A1(D[5]), .A2(n_0_16), .B1(n_0_15), .B2(Q[5]), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_6));
   AOI22_X1 i_0_13 (.A1(D[6]), .A2(n_0_16), .B1(n_0_15), .B2(Q[6]), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_7));
   AOI22_X1 i_0_15 (.A1(D[7]), .A2(n_0_16), .B1(n_0_15), .B2(Q[7]), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_8));
   AOI22_X1 i_0_17 (.A1(D[8]), .A2(n_0_16), .B1(n_0_15), .B2(Q[8]), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_9));
   AOI22_X1 i_0_19 (.A1(D[9]), .A2(n_0_16), .B1(n_0_15), .B2(Q[9]), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_10));
   AOI22_X1 i_0_21 (.A1(D[10]), .A2(n_0_16), .B1(n_0_15), .B2(Q[10]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_11));
   AOI22_X1 i_0_23 (.A1(D[11]), .A2(n_0_16), .B1(n_0_15), .B2(Q[11]), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_12));
   AOI22_X1 i_0_25 (.A1(D[12]), .A2(n_0_16), .B1(n_0_15), .B2(Q[12]), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_13));
   AOI22_X1 i_0_27 (.A1(D[13]), .A2(n_0_16), .B1(n_0_15), .B2(Q[13]), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_14));
   AOI22_X1 i_0_29 (.A1(D[14]), .A2(n_0_16), .B1(n_0_15), .B2(Q[14]), .ZN(n_0_14));
   NOR2_X1 i_0_30 (.A1(rst), .A2(load), .ZN(n_0_15));
   NOR2_X1 i_0_31 (.A1(n_0_17), .A2(rst), .ZN(n_0_16));
   INV_X1 i_0_32 (.A(load), .ZN(n_0_17));
   INV_X1 i_0_33 (.A(Clk), .ZN(n_15));
endmodule

module Euler(M1Data1, M2Data1, M1Data1W, M2Data1W, M1Data2, M2Data2, M1Address1, 
      M1Address2, M2Address1, M2Address2, Un, Uz, Ti, Uk, h_to_interpolation, 
      h_in, clk, rst, processCMD, Var1, Var2, Var3, Var4, Var5, selector, 
      Shift_Interpolation, writeX, writeU, programDone, Failure);
   input [63:0]M1Data1;
   input [63:0]M2Data1;
   output [63:0]M1Data1W;
   output [63:0]M2Data1W;
   input [63:0]M1Data2;
   input [63:0]M2Data2;
   output [15:0]M1Address1;
   output [15:0]M1Address2;
   output [15:0]M2Address1;
   output [15:0]M2Address2;
   output [15:0]Un;
   output [15:0]Uz;
   output [15:0]Ti;
   input [15:0]Uk;
   output [15:0]h_to_interpolation;
   input [15:0]h_in;
   input clk;
   input rst;
   input processCMD;
   input Var1;
   input Var2;
   input Var3;
   input Var4;
   input Var5;
   input [2:0]selector;
   output Shift_Interpolation;
   output writeX;
   output writeU;
   output programDone;
   output Failure;

   wire vectorDone;
   wire [15:0]Add_XpreS;
   wire doneB;
   wire [15:0]Add_B;
   wire firstRaw;
   wire doneA;
   wire [15:0]Add_A;
   wire [15:0]Add_xs1;
   wire [15:0]Add_xs2;
   wire [15:0]Add_X;
   wire [15:0]Add_XpreR;
   wire [15:0]Add_Ucalc;
   wire [15:0]Add_Un;
   wire [15:0]Add_Uz;
   wire overflow2;
   wire overflow1;
   wire VariableStep;
   wire n_0_0;
   wire n_0_1;
   wire decOut;
   wire [15:0]to_U;
   wire [15:0]B;
   wire [15:0]A;
   wire [15:0]Xn;
   wire resetA_B;
   wire elementDone;
   wire n_0_3_0;
   wire n_0_3_1;
   wire XstoreCounterEnable;
   wire n_0_3_2;
   wire XS1CounterEnable;
   wire n_0_3_3;
   wire XS2CounterEnable;
   wire incXR;
   wire U_enable;

   assign M1Data1W[63] = 1'b0;
   assign M1Data1W[62] = 1'b0;
   assign M1Data1W[61] = 1'b0;
   assign M1Data1W[60] = 1'b0;
   assign M1Data1W[59] = 1'b0;
   assign M1Data1W[58] = 1'b0;
   assign M1Data1W[57] = 1'b0;
   assign M1Data1W[56] = 1'b0;
   assign M1Data1W[55] = 1'b0;
   assign M1Data1W[54] = 1'b0;
   assign M1Data1W[53] = 1'b0;
   assign M1Data1W[52] = 1'b0;
   assign M1Data1W[51] = 1'b0;
   assign M1Data1W[50] = 1'b0;
   assign M1Data1W[49] = 1'b0;
   assign M1Data1W[48] = 1'b0;
   assign M1Data1W[47] = 1'b0;
   assign M1Data1W[46] = 1'b0;
   assign M1Data1W[45] = 1'b0;
   assign M1Data1W[44] = 1'b0;
   assign M1Data1W[43] = 1'b0;
   assign M1Data1W[42] = 1'b0;
   assign M1Data1W[41] = 1'b0;
   assign M1Data1W[40] = 1'b0;
   assign M1Data1W[39] = 1'b0;
   assign M1Data1W[38] = 1'b0;
   assign M1Data1W[37] = 1'b0;
   assign M1Data1W[36] = 1'b0;
   assign M1Data1W[35] = 1'b0;
   assign M1Data1W[34] = 1'b0;
   assign M1Data1W[33] = 1'b0;
   assign M1Data1W[32] = 1'b0;
   assign M1Data1W[31] = 1'b0;
   assign M1Data1W[30] = 1'b0;
   assign M1Data1W[29] = 1'b0;
   assign M1Data1W[28] = 1'b0;
   assign M1Data1W[27] = 1'b0;
   assign M1Data1W[26] = 1'b0;
   assign M1Data1W[25] = 1'b0;
   assign M1Data1W[24] = 1'b0;
   assign M1Data1W[23] = 1'b0;
   assign M1Data1W[22] = 1'b0;
   assign M1Data1W[21] = 1'b0;
   assign M1Data1W[20] = 1'b0;
   assign M1Data1W[19] = 1'b0;
   assign M1Data1W[18] = 1'b0;
   assign M1Data1W[17] = 1'b0;
   assign M1Data1W[16] = 1'b0;
   assign M2Data1W[63] = 1'b0;
   assign M2Data1W[62] = 1'b0;
   assign M2Data1W[61] = 1'b0;
   assign M2Data1W[60] = 1'b0;
   assign M2Data1W[59] = 1'b0;
   assign M2Data1W[58] = 1'b0;
   assign M2Data1W[57] = 1'b0;
   assign M2Data1W[56] = 1'b0;
   assign M2Data1W[55] = 1'b0;
   assign M2Data1W[54] = 1'b0;
   assign M2Data1W[53] = 1'b0;
   assign M2Data1W[52] = 1'b0;
   assign M2Data1W[51] = 1'b0;
   assign M2Data1W[50] = 1'b0;
   assign M2Data1W[49] = 1'b0;
   assign M2Data1W[48] = 1'b0;
   assign M2Data1W[47] = 1'b0;
   assign M2Data1W[46] = 1'b0;
   assign M2Data1W[45] = 1'b0;
   assign M2Data1W[44] = 1'b0;
   assign M2Data1W[43] = 1'b0;
   assign M2Data1W[42] = 1'b0;
   assign M2Data1W[41] = 1'b0;
   assign M2Data1W[40] = 1'b0;
   assign M2Data1W[39] = 1'b0;
   assign M2Data1W[38] = 1'b0;
   assign M2Data1W[37] = 1'b0;
   assign M2Data1W[36] = 1'b0;
   assign M2Data1W[35] = 1'b0;
   assign M2Data1W[34] = 1'b0;
   assign M2Data1W[33] = 1'b0;
   assign M2Data1W[32] = 1'b0;
   assign M2Data1W[31] = 1'b0;
   assign M2Data1W[30] = 1'b0;
   assign M2Data1W[29] = 1'b0;
   assign M2Data1W[28] = 1'b0;
   assign M2Data1W[27] = 1'b0;
   assign M2Data1W[26] = 1'b0;
   assign M2Data1W[25] = 1'b0;
   assign M2Data1W[24] = 1'b0;
   assign M2Data1W[23] = 1'b0;
   assign M2Data1W[22] = 1'b0;
   assign M2Data1W[21] = 1'b0;
   assign M2Data1W[20] = 1'b0;
   assign M2Data1W[19] = 1'b0;
   assign M2Data1W[18] = 1'b0;
   assign M2Data1W[17] = 1'b0;
   assign M2Data1W[16] = 1'b0;
   assign Un[15] = M2Data1[15];
   assign Un[14] = M2Data1[14];
   assign Un[13] = M2Data1[13];
   assign Un[12] = M2Data1[12];
   assign Un[11] = M2Data1[11];
   assign Un[10] = M2Data1[10];
   assign Un[9] = M2Data1[9];
   assign Un[8] = M2Data1[8];
   assign Un[7] = M2Data1[7];
   assign Un[6] = M2Data1[6];
   assign Un[5] = M2Data1[5];
   assign Un[4] = M2Data1[4];
   assign Un[3] = M2Data1[3];
   assign Un[2] = M2Data1[2];
   assign Un[1] = M2Data1[1];
   assign Un[0] = M2Data1[0];
   assign Uz[15] = M2Data2[15];
   assign Uz[14] = M2Data2[14];
   assign Uz[13] = M2Data2[13];
   assign Uz[12] = M2Data2[12];
   assign Uz[11] = M2Data2[11];
   assign Uz[10] = M2Data2[10];
   assign Uz[9] = M2Data2[9];
   assign Uz[8] = M2Data2[8];
   assign Uz[7] = M2Data2[7];
   assign Uz[6] = M2Data2[6];
   assign Uz[5] = M2Data2[5];
   assign Uz[4] = M2Data2[4];
   assign Uz[3] = M2Data2[3];
   assign Uz[2] = M2Data2[2];
   assign Uz[1] = M2Data2[1];
   assign Uz[0] = M2Data2[0];
   assign programDone = 1'b1;

   counter Xstore (.dataIn(), .offset({uc_0, uc_1, uc_2, n_5, n_4, n_3, n_2, n_1, 
      n_0, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9}), .load(), .enable(
      XstoreCounterEnable), .CLK(clk), .reset(), .universalReset(rst), .continue(), 
      .dataOut(Add_XpreS), .done(vectorDone), .NFN());
   counter__1_478 Bcounter (.dataIn(), .offset({uc_10, uc_11, uc_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18, uc_19}), 
      .load(), .enable(n_14), .CLK(clk), .reset(), .universalReset(resetA_B), 
      .continue(elementDone), .dataOut(Add_B), .done(doneB), .NFN());
   counter__14_425 Acounter (.dataIn(), .offset({uc_20, uc_21, uc_22, n_5, n_4, 
      n_3, n_2, n_1, n_0, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29}), 
      .load(), .enable(n_15), .CLK(clk), .reset(), .universalReset(resetA_B), 
      .continue(elementDone), .dataOut(Add_A), .done(doneA), .NFN(firstRaw));
   counter__16_425 XS1Counter (.dataIn(), .offset({uc_30, uc_31, uc_32, n_5, n_4, 
      n_3, n_2, n_1, n_0, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39}), 
      .load(), .enable(XS1CounterEnable), .CLK(clk), .reset(vectorDone), 
      .universalReset(rst), .continue(), .dataOut(Add_xs1), .done(), .NFN());
   counter__16_425__1 XS2Counter (.dataIn(), .offset({uc_40, uc_41, uc_42, n_5, 
      n_4, n_3, n_2, n_1, n_0, uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49}), 
      .load(), .enable(XS2CounterEnable), .CLK(clk), .reset(vectorDone), 
      .universalReset(rst), .continue(), .dataOut(Add_xs2), .done(), .NFN());
   counter__17_425 x (.dataIn(), .offset({uc_50, uc_51, uc_52, n_5, n_4, n_3, 
      n_2, n_1, n_0, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59}), .load(), 
      .enable(n_15), .CLK(clk), .reset(elementDone), .universalReset(rst), 
      .continue(), .dataOut(Add_X), .done(), .NFN());
   counter__18_425 XpreRead (.dataIn(), .offset({uc_60, uc_61, uc_62, n_5, n_4, 
      n_3, n_2, n_1, n_0, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69}), 
      .load(), .enable(incXR), .CLK(clk), .reset(), .universalReset(rst), 
      .continue(vectorDone), .dataOut(Add_XpreR), .done(), .NFN());
   counter__19_425 Ucalc (.dataIn(), .offset({uc_70, uc_71, uc_72, n_11, n_10, 
      n_9, n_8, n_7, n_6, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79}), 
      .load(), .enable(n_13), .CLK(clk), .reset(elementDone), .universalReset(
      rst), .continue(), .dataOut(Add_Ucalc), .done(), .NFN());
   counter__20_425 UnCounter (.dataIn(), .offset({uc_80, uc_81, uc_82, n_11, 
      n_10, n_9, n_8, n_7, n_6, uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89}), 
      .load(), .enable(n_12), .CLK(clk), .reset(elementDone), .universalReset(
      rst), .continue(), .dataOut(Add_Un), .done(), .NFN());
   counter__21_425 UZCounter (.dataIn(), .offset({uc_90, uc_91, uc_92, n_11, 
      n_10, n_9, n_8, n_7, n_6, uc_93, uc_94, uc_95, uc_96, uc_97, uc_98, uc_99}), 
      .load(), .enable(n_12), .CLK(clk), .reset(elementDone), .universalReset(
      rst), .continue(), .dataOut(Add_Uz), .done(), .NFN());
   booth_multiplier B_U_block (.m(B), .r({uc_100, M2Data1W[14], M2Data1W[13], 
      M2Data1W[12], M2Data1W[11], M2Data1W[10], M2Data1W[9], M2Data1W[8], 
      M2Data1W[7], M2Data1W[6], M2Data1W[5], M2Data1W[4], M2Data1W[3], 
      M2Data1W[2], M2Data1W[1], M2Data1W[0]}), .result(), .overflow(overflow2));
   booth_multiplier__1 A_X_block (.m(A), .r({uc_101, Xn[14], Xn[13], Xn[12], 
      Xn[11], Xn[10], Xn[9], Xn[8], Xn[7], Xn[6], Xn[5], Xn[4], Xn[3], Xn[2], 
      Xn[1], Xn[0]}), .result(), .overflow(overflow1));
   reg__3_24 Initreg (.D({uc_102, uc_103, uc_104, M1Data2[12], M1Data2[11], 
      M1Data2[10], M1Data2[9], M1Data2[8], M1Data2[7], M1Data2[6], M1Data2[5], 
      M1Data2[4], M1Data2[3], M1Data2[2], M1Data2[1], M1Data2[0]}), .load(decOut), 
      .Clk(clk), .Q({uc_105, uc_106, uc_107, VariableStep, n_11, n_10, n_9, n_8, 
      n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .rst(rst));
   Decoder1 busDec (.s(selector), .firstRaw(firstRaw), .d({decOut, uc_108, 
      uc_109, n_15, n_14, Shift_Interpolation, n_13, n_12, n_0_1, n_0_0}));
   reg__3_44 XprevReg (.D({M1Data2[15], M1Data2[14], M1Data2[13], M1Data2[12], 
      M1Data2[11], M1Data2[10], M1Data2[9], M1Data2[8], M1Data2[7], M1Data2[6], 
      M1Data2[5], M1Data2[4], M1Data2[3], M1Data2[2], M1Data2[1], M1Data2[0]}), 
      .load(n_0_1), .Clk(clk), .Q({M1Data1W[15], M1Data1W[14], M1Data1W[13], 
      M1Data1W[12], M1Data1W[11], M1Data1W[10], M1Data1W[9], M1Data1W[8], 
      M1Data1W[7], M1Data1W[6], M1Data1W[5], M1Data1W[4], M1Data1W[3], 
      M1Data1W[2], M1Data1W[1], M1Data1W[0]}), .rst(rst));
   twoInpMux UMux (.In0(Uk), .In1({M2Data1[15], M2Data1[14], M2Data1[13], 
      M2Data1[12], M2Data1[11], M2Data1[10], M2Data1[9], M2Data1[8], M2Data1[7], 
      M2Data1[6], M2Data1[5], M2Data1[4], M2Data1[3], M2Data1[2], M2Data1[1], 
      M2Data1[0]}), .selector(n_13), .out1(to_U));
   reg__3_64 Ureg (.D(to_U), .load(U_enable), .Clk(clk), .Q({M2Data1W[15], 
      M2Data1W[14], M2Data1W[13], M2Data1W[12], M2Data1W[11], M2Data1W[10], 
      M2Data1W[9], M2Data1W[8], M2Data1W[7], M2Data1W[6], M2Data1W[5], 
      M2Data1W[4], M2Data1W[3], M2Data1W[2], M2Data1W[1], M2Data1W[0]}), 
      .rst(rst));
   M1Add1Mux M1A1 (.Init(), .E(), .Ti(), .A(Add_A), .Xstore(Add_XpreS), .XS1(
      Add_xs1), .XS2(Add_xs2), .selector(selector), .Var1(Var1), .Var2(Var2), 
      .Var3(Var3), .Add(M1Address1));
   M1Add2Mux M1A2 (.H(), .Xn(Add_X), .Xprev(Add_XpreR), .Xs2(Add_xs2), .selector(
      selector), .Add(M1Address2));
   M2Add1Mux M2A1 (.Ucalc(Add_Ucalc), .Un(Add_Un), .Ustore(), .selector(selector), 
      .firstRaw(firstRaw), .Add(M2Address1));
   M2Add2Mux M2A2 (.B(Add_B), .Uz(Add_Uz), .selector(selector), .firstRaw(
      firstRaw), .Add(M2Address2));
   reg__3_84 Breg (.D({M2Data2[15], M2Data2[14], M2Data2[13], M2Data2[12], 
      M2Data2[11], M2Data2[10], M2Data2[9], M2Data2[8], M2Data2[7], M2Data2[6], 
      M2Data2[5], M2Data2[4], M2Data2[3], M2Data2[2], M2Data2[1], M2Data2[0]}), 
      .load(n_14), .Clk(clk), .Q(B), .rst(rst));
   reg__3_104 Areg (.D({M1Data1[15], M1Data1[14], M1Data1[13], M1Data1[12], 
      M1Data1[11], M1Data1[10], M1Data1[9], M1Data1[8], M1Data1[7], M1Data1[6], 
      M1Data1[5], M1Data1[4], M1Data1[3], M1Data1[2], M1Data1[1], M1Data1[0]}), 
      .load(n_15), .Clk(clk), .Q(A), .rst(rst));
   reg__3_124 Xnreg (.D({uc_110, M1Data2[14], M1Data2[13], M1Data2[12], 
      M1Data2[11], M1Data2[10], M1Data2[9], M1Data2[8], M1Data2[7], M1Data2[6], 
      M1Data2[5], M1Data2[4], M1Data2[3], M1Data2[2], M1Data2[1], M1Data2[0]}), 
      .load(n_15), .Clk(clk), .Q({uc_111, Xn[14], Xn[13], Xn[12], Xn[11], Xn[10], 
      Xn[9], Xn[8], Xn[7], Xn[6], Xn[5], Xn[4], Xn[3], Xn[2], Xn[1], Xn[0]}), 
      .rst(rst));
   OR2_X1 i_0_2_0 (.A1(rst), .A2(vectorDone), .ZN(resetA_B));
   AND2_X1 i_0_2_1 (.A1(doneA), .A2(doneB), .ZN(elementDone));
   INV_X1 i_0_3_0 (.A(n_0_1), .ZN(n_0_3_0));
   INV_X1 i_0_3_1 (.A(Var4), .ZN(n_0_3_1));
   AOI21_X1 i_0_3_2 (.A(n_0_3_0), .B1(n_0_3_1), .B2(VariableStep), .ZN(
      XstoreCounterEnable));
   AOI21_X1 i_0_3_3 (.A(n_0_0), .B1(n_0_1), .B2(Var1), .ZN(n_0_3_2));
   INV_X1 i_0_3_4 (.A(n_0_3_2), .ZN(XS1CounterEnable));
   AOI21_X1 i_0_3_5 (.A(n_0_0), .B1(n_0_1), .B2(Var2), .ZN(n_0_3_3));
   INV_X1 i_0_3_6 (.A(n_0_3_3), .ZN(XS2CounterEnable));
   OR2_X1 i_0_3_7 (.A1(decOut), .A2(n_0_1), .ZN(incXR));
   OR2_X1 i_0_0_0 (.A1(overflow1), .A2(overflow2), .ZN(Failure));
   OR2_X1 i_0_1_0 (.A1(n_13), .A2(n_12), .ZN(U_enable));
endmodule
