/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 10:54:45 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 450013737 */

module mux__0_5079(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5082(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5085(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5088(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5091(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5094(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5097(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5100(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5103(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5106(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5109(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5112(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5115(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux__0_5118(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   AND2_X1 i_0_0 (.A1(i2), .A2(sel), .ZN(Carry));
   XOR2_X1 i_0_1 (.A(i2), .B(sel), .Z(out1));
endmodule

module mux(sel, in1, in2, i1, i2, out1, Carry);
   input sel;
   input in1;
   input in2;
   input i1;
   input i2;
   output out1;
   output Carry;

   XOR2_X1 i_1_0 (.A(in1), .B(sel), .Z(out1));
endmodule

module Addition1(A, B, Cin, sum, Cout);
   input [15:0]A;
   input [15:0]B;
   input Cin;
   output [15:0]sum;
   output Cout;

   mux__0_5079 muxx_1_muxx_j (.sel(B[0]), .in1(), .in2(), .i1(), .i2(B[1]), 
      .out1(sum[1]), .Carry(n_0));
   mux__0_5082 muxx_2_muxx_j (.sel(n_0), .in1(), .in2(), .i1(), .i2(B[2]), 
      .out1(sum[2]), .Carry(n_1));
   mux__0_5085 muxx_3_muxx_j (.sel(n_1), .in1(), .in2(), .i1(), .i2(B[3]), 
      .out1(sum[3]), .Carry(n_2));
   mux__0_5088 muxx_4_muxx_j (.sel(n_2), .in1(), .in2(), .i1(), .i2(B[4]), 
      .out1(sum[4]), .Carry(n_3));
   mux__0_5091 muxx_5_muxx_j (.sel(n_3), .in1(), .in2(), .i1(), .i2(B[5]), 
      .out1(sum[5]), .Carry(n_4));
   mux__0_5094 muxx_6_muxx_j (.sel(n_4), .in1(), .in2(), .i1(), .i2(B[6]), 
      .out1(sum[6]), .Carry(n_5));
   mux__0_5097 muxx_7_muxx_j (.sel(n_5), .in1(), .in2(), .i1(), .i2(B[7]), 
      .out1(sum[7]), .Carry(n_6));
   mux__0_5100 muxx_8_muxx_j (.sel(n_6), .in1(), .in2(), .i1(), .i2(B[8]), 
      .out1(sum[8]), .Carry(n_7));
   mux__0_5103 muxx_9_muxx_j (.sel(n_7), .in1(), .in2(), .i1(), .i2(B[9]), 
      .out1(sum[9]), .Carry(n_8));
   mux__0_5106 muxx_10_muxx_j (.sel(n_8), .in1(), .in2(), .i1(), .i2(B[10]), 
      .out1(sum[10]), .Carry(n_9));
   mux__0_5109 muxx_11_muxx_j (.sel(n_9), .in1(), .in2(), .i1(), .i2(B[11]), 
      .out1(sum[11]), .Carry(n_10));
   mux__0_5112 muxx_12_muxx_j (.sel(n_10), .in1(), .in2(), .i1(), .i2(B[12]), 
      .out1(sum[12]), .Carry(n_11));
   mux__0_5115 muxx_13_muxx_j (.sel(n_11), .in1(), .in2(), .i1(), .i2(B[13]), 
      .out1(sum[13]), .Carry(n_12));
   mux__0_5118 muxx_14_muxx_j (.sel(n_12), .in1(), .in2(), .i1(), .i2(B[14]), 
      .out1(sum[14]), .Carry(n_13));
   mux muxx_15_muxx_j (.sel(n_13), .in1(B[15]), .in2(), .i1(), .i2(), .out1(
      sum[15]), .Carry());
endmodule

module Partial_Full_Adder__0_675(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_671(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_667(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_663(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_659(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_655(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_651(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_647(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_643(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_639(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_635(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_631(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_627(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_623(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_619(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_615(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_708(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_675 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_671 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_667 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_663 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_659 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_655 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_651 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_647 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_643 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_639 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_635 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_631 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_627 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_623 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_619 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_615 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_843(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_839(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_835(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_831(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_827(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_823(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_819(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_815(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_811(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_807(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_803(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_799(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_795(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_791(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_787(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_783(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_876(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_843 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_839 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_835 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_831 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_827 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_823 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_819 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_815 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_811 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_807 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_803 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_799 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_795 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_791 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_787 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_783 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_1011(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1007(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1003(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_999(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_995(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_991(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_987(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_983(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_979(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_975(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_971(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_967(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_963(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_959(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_955(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_951(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_1044(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_1011 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_1007 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_1003 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_999 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_995 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_991 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_987 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_983 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_979 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_975 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_971 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_967 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_963 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_959 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_955 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_951 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_1179(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1175(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1171(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1167(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1163(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1159(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1155(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1151(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1147(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1143(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1139(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1135(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1131(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1127(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1123(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1119(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_1212(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_1179 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_1175 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_1171 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1167 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1163 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1159 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1155 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1151 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1147 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1143 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1139 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1135 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1131 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1127 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1123 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1119 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_1347(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1343(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1339(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1335(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1331(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1327(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1323(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1319(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1315(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1311(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1307(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1303(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1299(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1295(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1291(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1287(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_1380(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_1347 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_1343 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_1339 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1335 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1331 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1327 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1323 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1319 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1315 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1311 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1307 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1303 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1299 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1295 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1291 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1287 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_1515(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1511(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1507(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1503(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1499(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1495(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1491(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1487(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1483(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1479(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1475(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1471(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1467(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1463(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1459(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1455(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_1548(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_1515 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_1511 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_1507 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1503 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1499 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1495 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1491 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1487 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1483 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1479 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1475 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1471 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1467 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1463 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1459 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1455 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_1683(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1679(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1675(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1671(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1667(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1663(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1659(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1655(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1651(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1647(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1643(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1639(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1635(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1631(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1627(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1623(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_1716(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_1683 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_1679 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_1675 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1671 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1667 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1663 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1659 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1655 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1651 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1647 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1643 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1639 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1635 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1631 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1627 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1623 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_1851(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1847(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1843(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1839(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1835(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1831(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1827(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1823(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1819(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1815(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1811(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1807(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1803(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1799(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1795(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1791(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_1884(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_1851 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_1847 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_1843 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1839 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1835 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1831 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1827 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1823 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1819 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1815 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1811 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1807 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1803 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1799 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1795 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1791 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_2019(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2015(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2011(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2007(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2003(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1999(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1995(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1991(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1987(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1983(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1979(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1975(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1971(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1967(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1963(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1959(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_2052(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_2019 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_2015 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_2011 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2007 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2003 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1999 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1995 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1991 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1987 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1983 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1979 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1975 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1971 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1967 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1963 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1959 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_2187(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2183(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2179(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2175(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2171(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2167(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2163(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2159(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2155(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2151(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2147(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2143(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2139(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2135(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2131(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2127(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_2220(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_2187 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_2183 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_2179 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2175 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2171 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2167 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2163 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2159 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2155 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2151 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2147 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2143 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2139 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2135 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2131 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2127 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_2355(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2351(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2347(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2343(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2339(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2335(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2331(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2327(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2323(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2319(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2315(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2311(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2307(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2303(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2299(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2295(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_2388(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_2355 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_2351 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_2347 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2343 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2339 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2335 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2331 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2327 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2323 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2319 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2315 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2311 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2307 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2303 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2299 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2295 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_2523(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2519(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2515(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2511(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2507(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2503(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2499(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2495(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2491(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2487(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2483(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2479(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2475(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2471(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2467(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2463(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   AND2_X1 i_2_0 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_2556(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_2523 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_2519 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_2515 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2511 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2507 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2503 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2499 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2495 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2491 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2487 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2483 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2479 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2475 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2471 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2467 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2463 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_2691(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2687(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2683(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2679(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2675(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2671(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2667(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2663(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2659(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2655(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2651(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2647(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2643(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2639(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2635(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2631(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_2724(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_2691 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_2687 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_2683 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2679 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2675 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2671 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2667 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2663 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2659 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2655 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2651 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2647 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2643 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2639 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2635 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2631 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_2859(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2855(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2851(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2847(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2843(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2839(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2835(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2831(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2827(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2823(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2819(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2815(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2811(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2807(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2803(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2799(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_2892(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_2859 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_2855 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_2851 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2847 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2843 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2839 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2835 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2831 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2827 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2823 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2819 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2815 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2811 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2807 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2803 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2799 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_3027(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_3023(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3019(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3015(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3011(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3007(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3003(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2999(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2995(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2991(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2987(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2983(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2979(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2975(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2971(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2967(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_3060(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_3027 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_3023 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_3019 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_3015 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_3011 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_3007 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_3003 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2999 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2995 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2991 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2987 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2983 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2979 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2975 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2971 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2967 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_3195(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_3191(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3187(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3183(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3179(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3175(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3171(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3167(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3163(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3159(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3155(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3151(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3147(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3143(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3139(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3135(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_3228(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_3195 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_3191 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_3187 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_3183 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_3179 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_3175 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_3171 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_3167 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_3163 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_3159 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_3155 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_3151 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_3147 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_3143 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_3139 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_3135 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_3363(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_3359(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3355(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3351(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3347(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3343(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3339(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3335(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3331(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3327(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3323(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3319(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3315(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3311(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3307(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3303(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_3396(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_3363 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_3359 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_3355 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_3351 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_3347 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_3343 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_3339 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_3335 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_3331 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_3327 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_3323 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_3319 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_3315 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_3311 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_3307 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_3303 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_3531(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_3527(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3523(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3519(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3515(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3511(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3507(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3503(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3499(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3495(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3491(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3487(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3483(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3479(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3475(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3471(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_3564(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_3531 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_3527 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_3523 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_3519 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_3515 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_3511 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_3507 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_3503 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_3499 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_3495 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_3491 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_3487 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_3483 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_3479 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_3475 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_3471 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_3699(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_3695(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3691(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3687(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3683(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3679(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3675(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3671(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3667(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3663(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3659(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3655(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3651(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3647(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3643(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3639(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_3732(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_3699 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_3695 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_3691 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_3687 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_3683 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_3679 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_3675 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_3671 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_3667 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_3663 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_3659 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_3655 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_3651 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_3647 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_3643 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_3639 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_3867(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_3863(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3859(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3855(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3851(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3847(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3843(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3839(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3835(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3831(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3827(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3823(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3819(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3815(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3811(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3807(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_3900(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_3867 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_3863 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_3859 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_3855 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_3851 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_3847 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_3843 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_3839 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_3835 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_3831 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_3827 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_3823 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_3819 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_3815 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_3811 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_3807 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_4035(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_4031(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4027(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4023(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4019(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4015(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4011(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4007(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4003(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3999(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3995(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3991(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3987(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3983(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3979(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_3975(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_4068(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_4035 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_4031 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_4027 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_4023 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_4019 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_4015 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_4011 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_4007 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_4003 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_3999 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_3995 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_3991 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_3987 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_3983 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_3979 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_3975 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_4203(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_4199(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4195(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4191(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4187(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4183(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4179(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4175(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4171(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4167(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4163(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4159(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4155(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4151(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4147(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4143(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_4236(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_4203 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_4199 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_4195 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_4191 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_4187 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_4183 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_4179 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_4175 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_4171 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_4167 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_4163 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_4159 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_4155 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_4151 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_4147 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_4143 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_4371(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_4367(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4363(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4359(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4355(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4351(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4347(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4343(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4339(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4335(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4331(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4327(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4323(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4319(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4315(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4311(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_4404(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_4371 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_4367 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_4363 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_4359 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_4355 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_4351 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_4347 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_4343 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_4339 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_4335 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_4331 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_4327 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_4323 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_4319 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_4315 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_4311 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_4539(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_4535(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4531(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4527(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4523(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4519(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4515(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4511(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4507(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4503(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4499(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4495(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4491(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4487(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4483(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4479(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_4572(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_4539 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_4535 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_4531 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_4527 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_4523 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_4519 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_4515 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_4511 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_4507 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_4503 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_4499 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_4495 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_4491 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_4487 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_4483 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_4479 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_4707(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_4703(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4699(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4695(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4691(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4687(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4683(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4679(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4675(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4671(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4667(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4663(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4659(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4655(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4651(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4647(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_4740(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_4707 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_4703 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_4699 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_4695 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_4691 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_4687 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_4683 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_4679 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_4675 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_4671 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_4667 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_4663 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_4659 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_4655 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_4651 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_4647 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_4875(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_4871(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4867(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4863(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4859(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4855(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4851(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4847(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4843(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4839(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4835(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4831(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4827(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4823(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4819(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4815(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_4908(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_4875 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_4871 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_4867 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_4863 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_4859 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_4855 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_4851 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_4847 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_4843 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_4839 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_4835 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_4831 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_4827 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_4823 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_4819 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_4815 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_5043(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_5039(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5035(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5031(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5027(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5023(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5019(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5015(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5011(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5007(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_5003(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4999(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4995(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4991(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4987(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_4983(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_5076(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_5043 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_5039 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_5035 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_5031 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_5027 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_5023 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_5019 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_5015 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_5011 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_5007 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_5003 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_4999 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_4995 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_4991 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_4987 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_4983 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module Partial_Full_Adder__0_80(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_84(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_88(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_92(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_96(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_100(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_104(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_108(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_112(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_116(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_120(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_124(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_128(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_132(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_136(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_140(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic(A, B, Cin, S, overFlow);
   input [32:0]A;
   input [32:0]B;
   input Cin;
   output [32:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire c;

   Partial_Full_Adder__0_80 GEN_FULL_ADDERS_32_FULL_ADDER_INST (.A(A[32]), 
      .B(B[32]), .Cin(c), .S(S[32]), .P(), .G());
   Partial_Full_Adder__0_84 GEN_FULL_ADDERS_31_FULL_ADDER_INST (.A(A[32]), 
      .B(B[31]), .Cin(n_39), .S(S[31]), .P(P), .G(G));
   Partial_Full_Adder__0_88 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_38), .S(S[30]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_92 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_37), .S(S[29]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_96 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_36), .S(S[28]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_100 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_35), .S(S[27]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_104 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_108 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_112 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_116 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_31), .S(S[23]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_120 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_30), .S(S[22]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_124 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_29), .S(S[21]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_128 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_28), .S(S[20]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_132 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_27), .S(S[19]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_136 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_26), .S(S[18]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_140 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(), .S(S[17]), .P(), .G(n_26));
   AOI21_X1 i_0_0 (.A(n_24), .B1(n_25), .B2(n_26), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(n_27));
   AOI21_X1 i_0_2 (.A(n_22), .B1(n_23), .B2(n_27), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_1), .ZN(n_28));
   AOI21_X1 i_0_4 (.A(n_20), .B1(n_21), .B2(n_28), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_29));
   AOI21_X1 i_0_6 (.A(n_18), .B1(n_19), .B2(n_29), .ZN(n_0_3));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_30));
   AOI21_X1 i_0_8 (.A(n_16), .B1(n_17), .B2(n_30), .ZN(n_0_4));
   INV_X1 i_0_9 (.A(n_0_4), .ZN(n_31));
   AOI21_X1 i_0_10 (.A(n_14), .B1(n_15), .B2(n_31), .ZN(n_0_5));
   INV_X1 i_0_11 (.A(n_0_5), .ZN(n_32));
   AOI21_X1 i_0_12 (.A(n_12), .B1(n_13), .B2(n_32), .ZN(n_0_6));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_33));
   AOI21_X1 i_0_14 (.A(n_10), .B1(n_11), .B2(n_33), .ZN(n_0_7));
   INV_X1 i_0_15 (.A(n_0_7), .ZN(n_34));
   AOI21_X1 i_0_16 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(n_0_8), .ZN(n_35));
   AOI21_X1 i_0_18 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_9), .ZN(n_36));
   AOI21_X1 i_0_20 (.A(n_4), .B1(n_5), .B2(n_36), .ZN(n_0_10));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_37));
   AOI21_X1 i_0_22 (.A(n_2), .B1(n_3), .B2(n_37), .ZN(n_0_11));
   INV_X1 i_0_23 (.A(n_0_11), .ZN(n_38));
   AOI21_X1 i_0_24 (.A(n_0), .B1(n_1), .B2(n_38), .ZN(n_0_12));
   INV_X1 i_0_25 (.A(n_0_12), .ZN(n_39));
   AOI21_X1 i_0_26 (.A(G), .B1(P), .B2(n_39), .ZN(n_0_13));
   INV_X1 i_0_27 (.A(n_0_13), .ZN(c));
endmodule

module booth_multiplier(m, r, result, overflow);
   input [15:0]m;
   input [15:0]r;
   output [15:0]result;
   output overflow;

   wire [15:0]mn;
   wire [32:0]\temp1[1] ;
   wire [32:0]\temp2[1] ;
   wire [32:0]\temp1[2] ;
   wire [32:0]\temp2[2] ;
   wire [32:0]\temp1[3] ;
   wire [32:0]\temp2[3] ;
   wire [32:0]\temp1[4] ;
   wire [32:0]\temp2[4] ;
   wire [32:0]\temp1[5] ;
   wire [32:0]\temp2[5] ;
   wire [32:0]\temp1[6] ;
   wire [32:0]\temp2[6] ;
   wire [32:0]\temp1[7] ;
   wire [32:0]\temp2[7] ;
   wire [32:0]\temp1[8] ;
   wire [32:0]\temp2[8] ;
   wire [32:0]\temp1[9] ;
   wire [32:0]\temp2[9] ;
   wire [32:0]\temp1[10] ;
   wire [32:0]\temp2[10] ;
   wire [32:0]\temp1[11] ;
   wire [32:0]\temp2[11] ;
   wire [32:0]\temp1[12] ;
   wire [32:0]\temp2[12] ;
   wire [32:0]\temp1[13] ;
   wire [32:0]\temp2[13] ;
   wire [32:0]\temp2[14] ;
   wire [32:0]\temp1[14] ;
   wire [15:0]notM;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_0;
   wire n_0_1_16;
   wire n_0_1;
   wire n_0_1_17;
   wire n_0_2;
   wire n_0_1_18;
   wire n_0_3;
   wire n_0_1_19;
   wire n_0_4;
   wire n_0_1_20;
   wire n_0_5;
   wire n_0_1_21;
   wire n_0_6;
   wire n_0_1_22;
   wire n_0_7;
   wire n_0_1_23;
   wire n_0_8;
   wire n_0_1_24;
   wire n_0_15;
   wire n_0_1_25;
   wire n_0_16;
   wire n_0_1_26;
   wire n_0_17;
   wire n_0_1_27;
   wire n_0_18;
   wire n_0_1_28;
   wire n_0_19;
   wire n_0_1_29;
   wire n_0_20;
   wire n_0_1_30;
   wire n_0_21;
   wire n_0_1_31;
   wire n_0_22;
   wire n_0_1_32;
   wire n_0_23;
   wire n_0_1_33;
   wire n_0_24;
   wire n_0_1_34;
   wire n_0_30;
   wire n_0_1_35;
   wire n_0_31;
   wire n_0_1_36;
   wire n_0_32;
   wire n_0_1_37;
   wire n_0_33;
   wire n_0_1_38;
   wire n_0_34;
   wire n_0_1_39;
   wire n_0_35;
   wire n_0_1_40;
   wire n_0_36;
   wire n_0_1_41;
   wire n_0_37;
   wire n_0_1_42;
   wire n_0_38;
   wire n_0_1_43;
   wire n_0_39;
   wire n_0_1_44;
   wire n_0_40;
   wire n_0_1_45;
   wire n_0_45;
   wire n_0_1_46;
   wire n_0_46;
   wire n_0_1_47;
   wire n_0_47;
   wire n_0_1_48;
   wire n_0_48;
   wire n_0_1_49;
   wire n_0_49;
   wire n_0_1_50;
   wire n_0_50;
   wire n_0_1_51;
   wire n_0_51;
   wire n_0_1_52;
   wire n_0_52;
   wire n_0_1_53;
   wire n_0_53;
   wire n_0_1_54;
   wire n_0_54;
   wire n_0_1_55;
   wire n_0_55;
   wire n_0_1_56;
   wire n_0_56;
   wire n_0_1_57;
   wire n_0_60;
   wire n_0_1_58;
   wire n_0_61;
   wire n_0_1_59;
   wire n_0_62;
   wire n_0_1_60;
   wire n_0_63;
   wire n_0_1_61;
   wire n_0_64;
   wire n_0_1_62;
   wire n_0_65;
   wire n_0_1_63;
   wire n_0_66;
   wire n_0_1_64;
   wire n_0_67;
   wire n_0_1_65;
   wire n_0_68;
   wire n_0_1_66;
   wire n_0_69;
   wire n_0_1_67;
   wire n_0_70;
   wire n_0_1_68;
   wire n_0_71;
   wire n_0_1_69;
   wire n_0_72;
   wire n_0_1_70;
   wire n_0_75;
   wire n_0_1_71;
   wire n_0_76;
   wire n_0_1_72;
   wire n_0_77;
   wire n_0_1_73;
   wire n_0_78;
   wire n_0_1_74;
   wire n_0_79;
   wire n_0_1_75;
   wire n_0_80;
   wire n_0_1_76;
   wire n_0_81;
   wire n_0_1_77;
   wire n_0_82;
   wire n_0_1_78;
   wire n_0_83;
   wire n_0_1_79;
   wire n_0_84;
   wire n_0_1_80;
   wire n_0_85;
   wire n_0_1_81;
   wire n_0_86;
   wire n_0_1_82;
   wire n_0_87;
   wire n_0_1_83;
   wire n_0_88;
   wire n_0_1_84;
   wire n_0_90;
   wire n_0_1_85;
   wire n_0_91;
   wire n_0_1_86;
   wire n_0_92;
   wire n_0_1_87;
   wire n_0_93;
   wire n_0_1_88;
   wire n_0_94;
   wire n_0_1_89;
   wire n_0_95;
   wire n_0_1_90;
   wire n_0_96;
   wire n_0_1_91;
   wire n_0_97;
   wire n_0_1_92;
   wire n_0_98;
   wire n_0_1_93;
   wire n_0_99;
   wire n_0_1_94;
   wire n_0_100;
   wire n_0_1_95;
   wire n_0_101;
   wire n_0_1_96;
   wire n_0_102;
   wire n_0_1_97;
   wire n_0_103;
   wire n_0_1_98;
   wire n_0_105;
   wire n_0_1_99;
   wire n_0_106;
   wire n_0_1_100;
   wire n_0_107;
   wire n_0_1_101;
   wire n_0_108;
   wire n_0_1_102;
   wire n_0_109;
   wire n_0_1_103;
   wire n_0_110;
   wire n_0_1_104;
   wire n_0_111;
   wire n_0_1_105;
   wire n_0_112;
   wire n_0_1_106;
   wire n_0_113;
   wire n_0_1_107;
   wire n_0_114;
   wire n_0_1_108;
   wire n_0_115;
   wire n_0_1_109;
   wire n_0_116;
   wire n_0_1_110;
   wire n_0_117;
   wire n_0_1_111;
   wire n_0_118;
   wire n_0_1_112;
   wire n_0_120;
   wire n_0_1_113;
   wire n_0_121;
   wire n_0_1_114;
   wire n_0_122;
   wire n_0_1_115;
   wire n_0_123;
   wire n_0_1_116;
   wire n_0_124;
   wire n_0_1_117;
   wire n_0_125;
   wire n_0_1_118;
   wire n_0_126;
   wire n_0_1_119;
   wire n_0_127;
   wire n_0_1_120;
   wire n_0_128;
   wire n_0_1_121;
   wire n_0_129;
   wire n_0_1_122;
   wire n_0_130;
   wire n_0_1_123;
   wire n_0_131;
   wire n_0_1_124;
   wire n_0_132;
   wire n_0_1_125;
   wire n_0_133;
   wire n_0_1_126;
   wire n_0_135;
   wire n_0_1_127;
   wire n_0_136;
   wire n_0_1_128;
   wire n_0_137;
   wire n_0_1_129;
   wire n_0_138;
   wire n_0_1_130;
   wire n_0_139;
   wire n_0_1_131;
   wire n_0_140;
   wire n_0_1_132;
   wire n_0_141;
   wire n_0_1_133;
   wire n_0_142;
   wire n_0_1_134;
   wire n_0_143;
   wire n_0_1_135;
   wire n_0_144;
   wire n_0_1_136;
   wire n_0_145;
   wire n_0_1_137;
   wire n_0_146;
   wire n_0_1_138;
   wire n_0_147;
   wire n_0_1_139;
   wire n_0_148;
   wire n_0_1_140;
   wire n_0_150;
   wire n_0_1_141;
   wire n_0_151;
   wire n_0_1_142;
   wire n_0_152;
   wire n_0_1_143;
   wire n_0_153;
   wire n_0_1_144;
   wire n_0_154;
   wire n_0_1_145;
   wire n_0_155;
   wire n_0_1_146;
   wire n_0_156;
   wire n_0_1_147;
   wire n_0_157;
   wire n_0_1_148;
   wire n_0_158;
   wire n_0_1_149;
   wire n_0_159;
   wire n_0_1_150;
   wire n_0_160;
   wire n_0_1_151;
   wire n_0_161;
   wire n_0_1_152;
   wire n_0_162;
   wire n_0_1_153;
   wire n_0_163;
   wire n_0_1_154;
   wire n_0_165;
   wire n_0_1_155;
   wire n_0_166;
   wire n_0_1_156;
   wire n_0_167;
   wire n_0_1_157;
   wire n_0_168;
   wire n_0_1_158;
   wire n_0_169;
   wire n_0_1_159;
   wire n_0_170;
   wire n_0_1_160;
   wire n_0_171;
   wire n_0_1_161;
   wire n_0_172;
   wire n_0_1_162;
   wire n_0_173;
   wire n_0_1_163;
   wire n_0_174;
   wire n_0_1_164;
   wire n_0_175;
   wire n_0_1_165;
   wire n_0_176;
   wire n_0_1_166;
   wire n_0_177;
   wire n_0_1_167;
   wire n_0_178;
   wire n_0_1_168;
   wire n_0_180;
   wire n_0_1_169;
   wire n_0_181;
   wire n_0_1_170;
   wire n_0_182;
   wire n_0_1_171;
   wire n_0_183;
   wire n_0_1_172;
   wire n_0_184;
   wire n_0_1_173;
   wire n_0_185;
   wire n_0_1_174;
   wire n_0_186;
   wire n_0_1_175;
   wire n_0_187;
   wire n_0_1_176;
   wire n_0_188;
   wire n_0_1_177;
   wire n_0_189;
   wire n_0_1_178;
   wire n_0_190;
   wire n_0_1_179;
   wire n_0_191;
   wire n_0_1_180;
   wire n_0_192;
   wire n_0_1_181;
   wire n_0_193;
   wire n_0_1_182;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_1_183;
   wire n_0_1_184;
   wire n_0_1_185;
   wire n_0_1_186;
   wire n_0_1_187;
   wire n_0_10;
   wire n_0_1_188;
   wire n_0_26;
   wire n_0_1_189;
   wire n_0_42;
   wire n_0_1_190;
   wire n_0_58;
   wire n_0_1_191;
   wire n_0_1_192;
   wire n_0_9;
   wire n_0_1_193;
   wire n_0_25;
   wire n_0_1_194;
   wire n_0_41;
   wire n_0_1_195;
   wire n_0_57;
   wire n_0_1_196;
   wire n_0_73;
   wire n_0_1_197;
   wire n_0_1_198;
   wire n_0_12;
   wire n_0_1_199;
   wire n_0_28;
   wire n_0_1_200;
   wire n_0_1_201;
   wire n_0_13;
   wire n_0_1_202;
   wire n_0_1_203;
   wire n_0_1_204;
   wire n_0_11;
   wire n_0_1_205;
   wire n_0_27;
   wire n_0_1_206;
   wire n_0_43;
   wire n_0_1_207;
   wire n_0_1_208;
   wire n_0_1_209;
   wire n_0_14;
   wire n_0_1_210;
   wire n_0_1_211;
   wire n_0_29;
   wire n_0_1_212;
   wire n_0_1_213;
   wire n_0_1_214;
   wire n_0_1_215;
   wire n_0_1_216;
   wire n_0_44;
   wire n_0_1_217;
   wire n_0_1_218;
   wire n_0_1_219;
   wire n_0_1_220;
   wire n_0_1_221;
   wire n_0_59;
   wire n_0_1_222;
   wire n_0_1_223;
   wire n_0_1_224;
   wire n_0_1_225;
   wire n_0_1_226;
   wire n_0_74;
   wire n_0_1_227;
   wire n_0_1_228;
   wire n_0_1_229;
   wire n_0_1_230;
   wire n_0_1_231;
   wire n_0_89;
   wire n_0_1_232;
   wire n_0_1_233;
   wire n_0_1_234;
   wire n_0_1_235;
   wire n_0_1_236;
   wire n_0_104;
   wire n_0_1_237;
   wire n_0_1_238;
   wire n_0_1_239;
   wire n_0_1_240;
   wire n_0_1_241;
   wire n_0_119;
   wire n_0_1_242;
   wire n_0_1_243;
   wire n_0_1_244;
   wire n_0_1_245;
   wire n_0_1_246;
   wire n_0_134;
   wire n_0_1_247;
   wire n_0_1_248;
   wire n_0_1_249;
   wire n_0_1_250;
   wire n_0_1_251;
   wire n_0_149;
   wire n_0_1_252;
   wire n_0_1_253;
   wire n_0_1_254;
   wire n_0_1_255;
   wire n_0_1_256;
   wire n_0_164;
   wire n_0_1_257;
   wire n_0_1_258;
   wire n_0_1_259;
   wire n_0_1_260;
   wire n_0_1_261;
   wire n_0_179;
   wire n_0_1_262;
   wire n_0_1_263;
   wire n_0_1_264;
   wire n_0_1_265;
   wire n_0_1_266;
   wire n_0_194;
   wire n_0_1_267;
   wire n_0_1_268;
   wire n_0_1_269;
   wire n_0_1_270;
   wire n_0_209;
   wire n_0_1_271;
   wire n_0_1_272;
   wire n_0_1_273;
   wire n_0_1_274;
   wire n_0_1_275;
   wire n_0_1_276;
   wire n_0_1_277;
   wire n_0_1_278;
   wire n_0_1_279;
   wire n_0_1_280;
   wire n_0_1_281;
   wire n_0_1_282;
   wire n_0_1_283;
   wire n_0_1_284;
   wire n_0_1_285;
   wire n_0_1_286;
   wire n_0_1_287;
   wire n_0_1_288;
   wire n_0_1_289;
   wire n_0_1_290;

   Addition1 U0 (.A(), .B(notM), .Cin(), .sum({mn[15], mn[14], mn[13], mn[12], 
      mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], 
      mn[1], uc_0}), .Cout());
   Carry_Look_Ahead_generic__0_708 x_1_Un (.A({n_0_209, uc_1, n_0_208, n_0_207, 
      n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, 
      n_0_198, n_0_197, n_0_196, n_0_195, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, uc_18}), 
      .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], m[7], m[6], m[5], 
      m[4], m[3], m[2], m[1], m[0], uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, 
      uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, 
      uc_35}), .Cin(), .S({\temp1[1] [32], \temp1[1] [31], \temp1[1] [30], 
      \temp1[1] [29], \temp1[1] [28], \temp1[1] [27], \temp1[1] [26], 
      \temp1[1] [25], \temp1[1] [24], \temp1[1] [23], \temp1[1] [22], 
      \temp1[1] [21], \temp1[1] [20], \temp1[1] [19], \temp1[1] [18], uc_36, 
      uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, 
      uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, uc_53}), .overFlow());
   Carry_Look_Ahead_generic__0_876 x_1_Ux (.A({n_0_209, uc_54, n_0_208, n_0_207, 
      n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, 
      n_0_198, n_0_197, n_0_196, n_0_195, uc_55, uc_56, uc_57, uc_58, uc_59, 
      uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, 
      uc_70, uc_71}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], mn[9], 
      mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], uc_72, uc_73, 
      uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, 
      uc_84, uc_85, uc_86, uc_87, uc_88}), .Cin(), .S({\temp2[1] [32], 
      \temp2[1] [31], \temp2[1] [30], \temp2[1] [29], \temp2[1] [28], 
      \temp2[1] [27], \temp2[1] [26], \temp2[1] [25], \temp2[1] [24], 
      \temp2[1] [23], \temp2[1] [22], \temp2[1] [21], \temp2[1] [20], 
      \temp2[1] [19], \temp2[1] [18], uc_89, uc_90, uc_91, uc_92, uc_93, uc_94, 
      uc_95, uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, 
      uc_105, uc_106}), .overFlow());
   Carry_Look_Ahead_generic__0_1044 x_2_Un (.A({n_0_194, uc_107, n_0_193, 
      n_0_192, n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, 
      n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, uc_108, uc_109, uc_110, 
      uc_111, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, uc_118, uc_119, 
      uc_120, uc_121, uc_122, uc_123, uc_124}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_125, uc_126, uc_127, uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, 
      uc_134, uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141}), .Cin(), 
      .S({\temp1[2] [32], \temp1[2] [31], \temp1[2] [30], \temp1[2] [29], 
      \temp1[2] [28], \temp1[2] [27], \temp1[2] [26], \temp1[2] [25], 
      \temp1[2] [24], \temp1[2] [23], \temp1[2] [22], \temp1[2] [21], 
      \temp1[2] [20], \temp1[2] [19], \temp1[2] [18], uc_142, uc_143, uc_144, 
      uc_145, uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, 
      uc_154, uc_155, uc_156, uc_157, uc_158, uc_159}), .overFlow());
   Carry_Look_Ahead_generic__0_1212 x_2_Ux (.A({n_0_194, uc_160, n_0_193, 
      n_0_192, n_0_191, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, 
      n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, uc_161, uc_162, uc_163, 
      uc_164, uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, uc_172, 
      uc_173, uc_174, uc_175, uc_176, uc_177}), .B({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], m[0], uc_178, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, 
      uc_185, uc_186, uc_187, uc_188, uc_189, uc_190, uc_191, uc_192, uc_193, 
      uc_194}), .Cin(), .S({\temp2[2] [32], \temp2[2] [31], \temp2[2] [30], 
      \temp2[2] [29], \temp2[2] [28], \temp2[2] [27], \temp2[2] [26], 
      \temp2[2] [25], \temp2[2] [24], \temp2[2] [23], \temp2[2] [22], 
      \temp2[2] [21], \temp2[2] [20], \temp2[2] [19], \temp2[2] [18], uc_195, 
      uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, uc_204, 
      uc_205, uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, uc_212}), 
      .overFlow());
   Carry_Look_Ahead_generic__0_1380 x_3_Un (.A({n_0_179, uc_213, n_0_178, 
      n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, 
      n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, uc_214, uc_215, uc_216, 
      uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, uc_223, uc_224, uc_225, 
      uc_226, uc_227, uc_228, uc_229, uc_230}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_231, uc_232, uc_233, uc_234, uc_235, uc_236, uc_237, uc_238, uc_239, 
      uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, uc_247}), .Cin(), 
      .S({\temp1[3] [32], \temp1[3] [31], \temp1[3] [30], \temp1[3] [29], 
      \temp1[3] [28], \temp1[3] [27], \temp1[3] [26], \temp1[3] [25], 
      \temp1[3] [24], \temp1[3] [23], \temp1[3] [22], \temp1[3] [21], 
      \temp1[3] [20], \temp1[3] [19], \temp1[3] [18], uc_248, uc_249, uc_250, 
      uc_251, uc_252, uc_253, uc_254, uc_255, uc_256, uc_257, uc_258, uc_259, 
      uc_260, uc_261, uc_262, uc_263, uc_264, uc_265}), .overFlow());
   Carry_Look_Ahead_generic__0_1548 x_3_Ux (.A({n_0_179, uc_266, n_0_178, 
      n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, 
      n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, uc_267, uc_268, uc_269, 
      uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, uc_278, 
      uc_279, uc_280, uc_281, uc_282, uc_283}), .B({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], m[0], uc_284, uc_285, uc_286, uc_287, uc_288, uc_289, uc_290, 
      uc_291, uc_292, uc_293, uc_294, uc_295, uc_296, uc_297, uc_298, uc_299, 
      uc_300}), .Cin(), .S({\temp2[3] [32], \temp2[3] [31], \temp2[3] [30], 
      \temp2[3] [29], \temp2[3] [28], \temp2[3] [27], \temp2[3] [26], 
      \temp2[3] [25], \temp2[3] [24], \temp2[3] [23], \temp2[3] [22], 
      \temp2[3] [21], \temp2[3] [20], \temp2[3] [19], \temp2[3] [18], uc_301, 
      uc_302, uc_303, uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, uc_310, 
      uc_311, uc_312, uc_313, uc_314, uc_315, uc_316, uc_317, uc_318}), 
      .overFlow());
   Carry_Look_Ahead_generic__0_1716 x_4_Un (.A({n_0_164, uc_319, n_0_163, 
      n_0_162, n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, 
      n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, uc_320, uc_321, uc_322, 
      uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, 
      uc_332, uc_333, uc_334, uc_335, uc_336}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_337, uc_338, uc_339, uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, 
      uc_346, uc_347, uc_348, uc_349, uc_350, uc_351, uc_352, uc_353}), .Cin(), 
      .S({\temp1[4] [32], \temp1[4] [31], \temp1[4] [30], \temp1[4] [29], 
      \temp1[4] [28], \temp1[4] [27], \temp1[4] [26], \temp1[4] [25], 
      \temp1[4] [24], \temp1[4] [23], \temp1[4] [22], \temp1[4] [21], 
      \temp1[4] [20], \temp1[4] [19], \temp1[4] [18], uc_354, uc_355, uc_356, 
      uc_357, uc_358, uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, 
      uc_366, uc_367, uc_368, uc_369, uc_370, uc_371}), .overFlow());
   Carry_Look_Ahead_generic__0_1884 x_4_Ux (.A({n_0_164, uc_372, n_0_163, 
      n_0_162, n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, 
      n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, uc_373, uc_374, uc_375, 
      uc_376, uc_377, uc_378, uc_379, uc_380, uc_381, uc_382, uc_383, uc_384, 
      uc_385, uc_386, uc_387, uc_388, uc_389}), .B({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], m[0], uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, 
      uc_397, uc_398, uc_399, uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, 
      uc_406}), .Cin(), .S({\temp2[4] [32], \temp2[4] [31], \temp2[4] [30], 
      \temp2[4] [29], \temp2[4] [28], \temp2[4] [27], \temp2[4] [26], 
      \temp2[4] [25], \temp2[4] [24], \temp2[4] [23], \temp2[4] [22], 
      \temp2[4] [21], \temp2[4] [20], \temp2[4] [19], \temp2[4] [18], uc_407, 
      uc_408, uc_409, uc_410, uc_411, uc_412, uc_413, uc_414, uc_415, uc_416, 
      uc_417, uc_418, uc_419, uc_420, uc_421, uc_422, uc_423, uc_424}), 
      .overFlow());
   Carry_Look_Ahead_generic__0_2052 x_5_Un (.A({n_0_149, uc_425, n_0_148, 
      n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, 
      n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, uc_426, uc_427, uc_428, 
      uc_429, uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, uc_436, uc_437, 
      uc_438, uc_439, uc_440, uc_441, uc_442}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, uc_450, uc_451, 
      uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, uc_459}), .Cin(), 
      .S({\temp1[5] [32], \temp1[5] [31], \temp1[5] [30], \temp1[5] [29], 
      \temp1[5] [28], \temp1[5] [27], \temp1[5] [26], \temp1[5] [25], 
      \temp1[5] [24], \temp1[5] [23], \temp1[5] [22], \temp1[5] [21], 
      \temp1[5] [20], \temp1[5] [19], \temp1[5] [18], uc_460, uc_461, uc_462, 
      uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, uc_469, uc_470, uc_471, 
      uc_472, uc_473, uc_474, uc_475, uc_476, uc_477}), .overFlow());
   Carry_Look_Ahead_generic__0_2220 x_5_Ux (.A({n_0_149, uc_478, n_0_148, 
      n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, 
      n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, uc_479, uc_480, uc_481, 
      uc_482, uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, 
      uc_491, uc_492, uc_493, uc_494, uc_495}), .B({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], m[0], uc_496, uc_497, uc_498, uc_499, uc_500, uc_501, uc_502, 
      uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, uc_509, uc_510, uc_511, 
      uc_512}), .Cin(), .S({\temp2[5] [32], \temp2[5] [31], \temp2[5] [30], 
      \temp2[5] [29], \temp2[5] [28], \temp2[5] [27], \temp2[5] [26], 
      \temp2[5] [25], \temp2[5] [24], \temp2[5] [23], \temp2[5] [22], 
      \temp2[5] [21], \temp2[5] [20], \temp2[5] [19], \temp2[5] [18], uc_513, 
      uc_514, uc_515, uc_516, uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, 
      uc_523, uc_524, uc_525, uc_526, uc_527, uc_528, uc_529, uc_530}), 
      .overFlow());
   Carry_Look_Ahead_generic__0_2388 x_6_Un (.A({n_0_134, uc_531, n_0_133, 
      n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, 
      n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, uc_532, uc_533, uc_534, 
      uc_535, uc_536, uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, 
      uc_544, uc_545, uc_546, uc_547, uc_548}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, uc_555, uc_556, uc_557, 
      uc_558, uc_559, uc_560, uc_561, uc_562, uc_563, uc_564, uc_565}), .Cin(), 
      .S({\temp1[6] [32], \temp1[6] [31], \temp1[6] [30], \temp1[6] [29], 
      \temp1[6] [28], \temp1[6] [27], \temp1[6] [26], \temp1[6] [25], 
      \temp1[6] [24], \temp1[6] [23], \temp1[6] [22], \temp1[6] [21], 
      \temp1[6] [20], \temp1[6] [19], \temp1[6] [18], uc_566, uc_567, uc_568, 
      uc_569, uc_570, uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, uc_577, 
      uc_578, uc_579, uc_580, uc_581, uc_582, uc_583}), .overFlow());
   Carry_Look_Ahead_generic__0_2556 x_6_Ux (.A({n_0_134, uc_584, n_0_133, 
      n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, 
      n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, uc_585, uc_586, uc_587, 
      uc_588, uc_589, uc_590, uc_591, uc_592, uc_593, uc_594, uc_595, uc_596, 
      uc_597, uc_598, uc_599, uc_600, uc_601}), .B({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], m[0], uc_602, uc_603, uc_604, uc_605, uc_606, uc_607, uc_608, 
      uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, uc_616, uc_617, 
      uc_618}), .Cin(), .S({\temp2[6] [32], \temp2[6] [31], \temp2[6] [30], 
      \temp2[6] [29], \temp2[6] [28], \temp2[6] [27], \temp2[6] [26], 
      \temp2[6] [25], \temp2[6] [24], \temp2[6] [23], \temp2[6] [22], 
      \temp2[6] [21], \temp2[6] [20], \temp2[6] [19], \temp2[6] [18], uc_619, 
      uc_620, uc_621, uc_622, uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, 
      uc_629, uc_630, uc_631, uc_632, uc_633, uc_634, uc_635, uc_636}), 
      .overFlow());
   Carry_Look_Ahead_generic__0_2724 x_7_Un (.A({n_0_119, uc_637, n_0_118, 
      n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
      n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, uc_638, uc_639, uc_640, 
      uc_641, uc_642, uc_643, uc_644, uc_645, uc_646, uc_647, uc_648, uc_649, 
      uc_650, uc_651, uc_652, uc_653, uc_654}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_655, uc_656, uc_657, uc_658, uc_659, uc_660, uc_661, uc_662, uc_663, 
      uc_664, uc_665, uc_666, uc_667, uc_668, uc_669, uc_670, uc_671}), .Cin(), 
      .S({\temp1[7] [32], \temp1[7] [31], \temp1[7] [30], \temp1[7] [29], 
      \temp1[7] [28], \temp1[7] [27], \temp1[7] [26], \temp1[7] [25], 
      \temp1[7] [24], \temp1[7] [23], \temp1[7] [22], \temp1[7] [21], 
      \temp1[7] [20], \temp1[7] [19], \temp1[7] [18], \temp1[7] [17], uc_672, 
      uc_673, uc_674, uc_675, uc_676, uc_677, uc_678, uc_679, uc_680, uc_681, 
      uc_682, uc_683, uc_684, uc_685, uc_686, uc_687, uc_688}), .overFlow());
   Carry_Look_Ahead_generic__0_2892 x_7_Ux (.A({n_0_119, uc_689, n_0_118, 
      n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, 
      n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, uc_690, uc_691, uc_692, 
      uc_693, uc_694, uc_695, uc_696, uc_697, uc_698, uc_699, uc_700, uc_701, 
      uc_702, uc_703, uc_704, uc_705, uc_706}), .B({mn[15], mn[14], mn[13], 
      mn[12], mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], 
      mn[2], mn[1], m[0], uc_707, uc_708, uc_709, uc_710, uc_711, uc_712, uc_713, 
      uc_714, uc_715, uc_716, uc_717, uc_718, uc_719, uc_720, uc_721, uc_722, 
      uc_723}), .Cin(), .S({\temp2[7] [32], \temp2[7] [31], \temp2[7] [30], 
      \temp2[7] [29], \temp2[7] [28], \temp2[7] [27], \temp2[7] [26], 
      \temp2[7] [25], \temp2[7] [24], \temp2[7] [23], \temp2[7] [22], 
      \temp2[7] [21], \temp2[7] [20], \temp2[7] [19], \temp2[7] [18], 
      \temp2[7] [17], uc_724, uc_725, uc_726, uc_727, uc_728, uc_729, uc_730, 
      uc_731, uc_732, uc_733, uc_734, uc_735, uc_736, uc_737, uc_738, uc_739, 
      uc_740}), .overFlow());
   Carry_Look_Ahead_generic__0_3060 x_8_Un (.A({n_0_104, uc_741, n_0_103, 
      n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, 
      n_0_93, n_0_92, n_0_91, n_0_90, uc_742, uc_743, uc_744, uc_745, uc_746, 
      uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, uc_753, uc_754, uc_755, 
      uc_756, uc_757, uc_758}), .B({m[15], m[14], m[13], m[12], m[11], m[10], 
      m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_759, uc_760, 
      uc_761, uc_762, uc_763, uc_764, uc_765, uc_766, uc_767, uc_768, uc_769, 
      uc_770, uc_771, uc_772, uc_773, uc_774, uc_775}), .Cin(), .S({
      \temp1[8] [32], \temp1[8] [31], \temp1[8] [30], \temp1[8] [29], 
      \temp1[8] [28], \temp1[8] [27], \temp1[8] [26], \temp1[8] [25], 
      \temp1[8] [24], \temp1[8] [23], \temp1[8] [22], \temp1[8] [21], 
      \temp1[8] [20], \temp1[8] [19], \temp1[8] [18], \temp1[8] [17], uc_776, 
      uc_777, uc_778, uc_779, uc_780, uc_781, uc_782, uc_783, uc_784, uc_785, 
      uc_786, uc_787, uc_788, uc_789, uc_790, uc_791, uc_792}), .overFlow());
   Carry_Look_Ahead_generic__0_3228 x_8_Ux (.A({n_0_104, uc_793, n_0_103, 
      n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, 
      n_0_93, n_0_92, n_0_91, n_0_90, uc_794, uc_795, uc_796, uc_797, uc_798, 
      uc_799, uc_800, uc_801, uc_802, uc_803, uc_804, uc_805, uc_806, uc_807, 
      uc_808, uc_809, uc_810}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], 
      mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], 
      m[0], uc_811, uc_812, uc_813, uc_814, uc_815, uc_816, uc_817, uc_818, 
      uc_819, uc_820, uc_821, uc_822, uc_823, uc_824, uc_825, uc_826, uc_827}), 
      .Cin(), .S({\temp2[8] [32], \temp2[8] [31], \temp2[8] [30], \temp2[8] [29], 
      \temp2[8] [28], \temp2[8] [27], \temp2[8] [26], \temp2[8] [25], 
      \temp2[8] [24], \temp2[8] [23], \temp2[8] [22], \temp2[8] [21], 
      \temp2[8] [20], \temp2[8] [19], \temp2[8] [18], \temp2[8] [17], uc_828, 
      uc_829, uc_830, uc_831, uc_832, uc_833, uc_834, uc_835, uc_836, uc_837, 
      uc_838, uc_839, uc_840, uc_841, uc_842, uc_843, uc_844}), .overFlow());
   Carry_Look_Ahead_generic__0_3396 x_9_Un (.A({n_0_89, uc_845, n_0_88, n_0_87, 
      n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, 
      n_0_77, n_0_76, n_0_75, uc_846, uc_847, uc_848, uc_849, uc_850, uc_851, 
      uc_852, uc_853, uc_854, uc_855, uc_856, uc_857, uc_858, uc_859, uc_860, 
      uc_861, uc_862}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], 
      m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_863, uc_864, uc_865, 
      uc_866, uc_867, uc_868, uc_869, uc_870, uc_871, uc_872, uc_873, uc_874, 
      uc_875, uc_876, uc_877, uc_878, uc_879}), .Cin(), .S({\temp1[9] [32], 
      \temp1[9] [31], \temp1[9] [30], \temp1[9] [29], \temp1[9] [28], 
      \temp1[9] [27], \temp1[9] [26], \temp1[9] [25], \temp1[9] [24], 
      \temp1[9] [23], \temp1[9] [22], \temp1[9] [21], \temp1[9] [20], 
      \temp1[9] [19], \temp1[9] [18], \temp1[9] [17], uc_880, uc_881, uc_882, 
      uc_883, uc_884, uc_885, uc_886, uc_887, uc_888, uc_889, uc_890, uc_891, 
      uc_892, uc_893, uc_894, uc_895, uc_896}), .overFlow());
   Carry_Look_Ahead_generic__0_3564 x_9_Ux (.A({n_0_89, uc_897, n_0_88, n_0_87, 
      n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, 
      n_0_77, n_0_76, n_0_75, uc_898, uc_899, uc_900, uc_901, uc_902, uc_903, 
      uc_904, uc_905, uc_906, uc_907, uc_908, uc_909, uc_910, uc_911, uc_912, 
      uc_913, uc_914}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], mn[10], 
      mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], m[0], 
      uc_915, uc_916, uc_917, uc_918, uc_919, uc_920, uc_921, uc_922, uc_923, 
      uc_924, uc_925, uc_926, uc_927, uc_928, uc_929, uc_930, uc_931}), .Cin(), 
      .S({\temp2[9] [32], \temp2[9] [31], \temp2[9] [30], \temp2[9] [29], 
      \temp2[9] [28], \temp2[9] [27], \temp2[9] [26], \temp2[9] [25], 
      \temp2[9] [24], \temp2[9] [23], \temp2[9] [22], \temp2[9] [21], 
      \temp2[9] [20], \temp2[9] [19], \temp2[9] [18], \temp2[9] [17], uc_932, 
      uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, uc_939, uc_940, uc_941, 
      uc_942, uc_943, uc_944, uc_945, uc_946, uc_947, uc_948}), .overFlow());
   Carry_Look_Ahead_generic__0_3732 x_10_Un (.A({n_0_74, uc_949, n_0_73, n_0_72, 
      n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, 
      n_0_62, n_0_61, n_0_60, uc_950, uc_951, uc_952, uc_953, uc_954, uc_955, 
      uc_956, uc_957, uc_958, uc_959, uc_960, uc_961, uc_962, uc_963, uc_964, 
      uc_965, uc_966}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], m[8], 
      m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_967, uc_968, uc_969, 
      uc_970, uc_971, uc_972, uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, 
      uc_979, uc_980, uc_981, uc_982, uc_983}), .Cin(), .S({\temp1[10] [32], 
      \temp1[10] [31], \temp1[10] [30], \temp1[10] [29], \temp1[10] [28], 
      \temp1[10] [27], \temp1[10] [26], \temp1[10] [25], \temp1[10] [24], 
      \temp1[10] [23], \temp1[10] [22], \temp1[10] [21], \temp1[10] [20], 
      \temp1[10] [19], \temp1[10] [18], \temp1[10] [17], uc_984, uc_985, uc_986, 
      uc_987, uc_988, uc_989, uc_990, uc_991, uc_992, uc_993, uc_994, uc_995, 
      uc_996, uc_997, uc_998, uc_999, uc_1000}), .overFlow());
   Carry_Look_Ahead_generic__0_3900 x_10_Ux (.A({n_0_74, uc_1001, n_0_73, n_0_72, 
      n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, 
      n_0_62, n_0_61, n_0_60, uc_1002, uc_1003, uc_1004, uc_1005, uc_1006, 
      uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, uc_1013, uc_1014, 
      uc_1015, uc_1016, uc_1017, uc_1018}), .B({mn[15], mn[14], mn[13], mn[12], 
      mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], 
      mn[1], m[0], uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, uc_1024, uc_1025, 
      uc_1026, uc_1027, uc_1028, uc_1029, uc_1030, uc_1031, uc_1032, uc_1033, 
      uc_1034, uc_1035}), .Cin(), .S({\temp2[10] [32], \temp2[10] [31], 
      \temp2[10] [30], \temp2[10] [29], \temp2[10] [28], \temp2[10] [27], 
      \temp2[10] [26], \temp2[10] [25], \temp2[10] [24], \temp2[10] [23], 
      \temp2[10] [22], \temp2[10] [21], \temp2[10] [20], \temp2[10] [19], 
      \temp2[10] [18], \temp2[10] [17], uc_1036, uc_1037, uc_1038, uc_1039, 
      uc_1040, uc_1041, uc_1042, uc_1043, uc_1044, uc_1045, uc_1046, uc_1047, 
      uc_1048, uc_1049, uc_1050, uc_1051, uc_1052}), .overFlow());
   Carry_Look_Ahead_generic__0_4068 x_11_Un (.A({n_0_59, uc_1053, n_0_58, n_0_57, 
      n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, 
      n_0_47, n_0_46, n_0_45, uc_1054, uc_1055, uc_1056, uc_1057, uc_1058, 
      uc_1059, uc_1060, uc_1061, uc_1062, uc_1063, uc_1064, uc_1065, uc_1066, 
      uc_1067, uc_1068, uc_1069, uc_1070}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_1071, uc_1072, uc_1073, uc_1074, uc_1075, uc_1076, uc_1077, uc_1078, 
      uc_1079, uc_1080, uc_1081, uc_1082, uc_1083, uc_1084, uc_1085, uc_1086, 
      uc_1087}), .Cin(), .S({\temp1[11] [32], \temp1[11] [31], \temp1[11] [30], 
      \temp1[11] [29], \temp1[11] [28], \temp1[11] [27], \temp1[11] [26], 
      \temp1[11] [25], \temp1[11] [24], \temp1[11] [23], \temp1[11] [22], 
      \temp1[11] [21], \temp1[11] [20], \temp1[11] [19], \temp1[11] [18], 
      \temp1[11] [17], uc_1088, uc_1089, uc_1090, uc_1091, uc_1092, uc_1093, 
      uc_1094, uc_1095, uc_1096, uc_1097, uc_1098, uc_1099, uc_1100, uc_1101, 
      uc_1102, uc_1103, uc_1104}), .overFlow());
   Carry_Look_Ahead_generic__0_4236 x_11_Ux (.A({n_0_59, uc_1105, n_0_58, n_0_57, 
      n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, 
      n_0_47, n_0_46, n_0_45, uc_1106, uc_1107, uc_1108, uc_1109, uc_1110, 
      uc_1111, uc_1112, uc_1113, uc_1114, uc_1115, uc_1116, uc_1117, uc_1118, 
      uc_1119, uc_1120, uc_1121, uc_1122}), .B({mn[15], mn[14], mn[13], mn[12], 
      mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], 
      mn[1], m[0], uc_1123, uc_1124, uc_1125, uc_1126, uc_1127, uc_1128, uc_1129, 
      uc_1130, uc_1131, uc_1132, uc_1133, uc_1134, uc_1135, uc_1136, uc_1137, 
      uc_1138, uc_1139}), .Cin(), .S({\temp2[11] [32], \temp2[11] [31], 
      \temp2[11] [30], \temp2[11] [29], \temp2[11] [28], \temp2[11] [27], 
      \temp2[11] [26], \temp2[11] [25], \temp2[11] [24], \temp2[11] [23], 
      \temp2[11] [22], \temp2[11] [21], \temp2[11] [20], \temp2[11] [19], 
      \temp2[11] [18], \temp2[11] [17], uc_1140, uc_1141, uc_1142, uc_1143, 
      uc_1144, uc_1145, uc_1146, uc_1147, uc_1148, uc_1149, uc_1150, uc_1151, 
      uc_1152, uc_1153, uc_1154, uc_1155, uc_1156}), .overFlow());
   Carry_Look_Ahead_generic__0_4404 x_12_Un (.A({n_0_44, uc_1157, n_0_43, n_0_42, 
      n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, 
      n_0_32, n_0_31, n_0_30, uc_1158, uc_1159, uc_1160, uc_1161, uc_1162, 
      uc_1163, uc_1164, uc_1165, uc_1166, uc_1167, uc_1168, uc_1169, uc_1170, 
      uc_1171, uc_1172, uc_1173, uc_1174}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_1175, uc_1176, uc_1177, uc_1178, uc_1179, uc_1180, uc_1181, uc_1182, 
      uc_1183, uc_1184, uc_1185, uc_1186, uc_1187, uc_1188, uc_1189, uc_1190, 
      uc_1191}), .Cin(), .S({\temp1[12] [32], \temp1[12] [31], \temp1[12] [30], 
      \temp1[12] [29], \temp1[12] [28], \temp1[12] [27], \temp1[12] [26], 
      \temp1[12] [25], \temp1[12] [24], \temp1[12] [23], \temp1[12] [22], 
      \temp1[12] [21], \temp1[12] [20], \temp1[12] [19], \temp1[12] [18], 
      \temp1[12] [17], uc_1192, uc_1193, uc_1194, uc_1195, uc_1196, uc_1197, 
      uc_1198, uc_1199, uc_1200, uc_1201, uc_1202, uc_1203, uc_1204, uc_1205, 
      uc_1206, uc_1207, uc_1208}), .overFlow());
   Carry_Look_Ahead_generic__0_4572 x_12_Ux (.A({n_0_44, uc_1209, n_0_43, n_0_42, 
      n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, 
      n_0_32, n_0_31, n_0_30, uc_1210, uc_1211, uc_1212, uc_1213, uc_1214, 
      uc_1215, uc_1216, uc_1217, uc_1218, uc_1219, uc_1220, uc_1221, uc_1222, 
      uc_1223, uc_1224, uc_1225, uc_1226}), .B({mn[15], mn[14], mn[13], mn[12], 
      mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], 
      mn[1], m[0], uc_1227, uc_1228, uc_1229, uc_1230, uc_1231, uc_1232, uc_1233, 
      uc_1234, uc_1235, uc_1236, uc_1237, uc_1238, uc_1239, uc_1240, uc_1241, 
      uc_1242, uc_1243}), .Cin(), .S({\temp2[12] [32], \temp2[12] [31], 
      \temp2[12] [30], \temp2[12] [29], \temp2[12] [28], \temp2[12] [27], 
      \temp2[12] [26], \temp2[12] [25], \temp2[12] [24], \temp2[12] [23], 
      \temp2[12] [22], \temp2[12] [21], \temp2[12] [20], \temp2[12] [19], 
      \temp2[12] [18], \temp2[12] [17], uc_1244, uc_1245, uc_1246, uc_1247, 
      uc_1248, uc_1249, uc_1250, uc_1251, uc_1252, uc_1253, uc_1254, uc_1255, 
      uc_1256, uc_1257, uc_1258, uc_1259, uc_1260}), .overFlow());
   Carry_Look_Ahead_generic__0_4740 x_13_Un (.A({n_0_29, uc_1261, n_0_28, n_0_27, 
      n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, uc_1262, uc_1263, uc_1264, uc_1265, uc_1266, 
      uc_1267, uc_1268, uc_1269, uc_1270, uc_1271, uc_1272, uc_1273, uc_1274, 
      uc_1275, uc_1276, uc_1277, uc_1278}), .B({m[15], m[14], m[13], m[12], 
      m[11], m[10], m[9], m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], 
      uc_1279, uc_1280, uc_1281, uc_1282, uc_1283, uc_1284, uc_1285, uc_1286, 
      uc_1287, uc_1288, uc_1289, uc_1290, uc_1291, uc_1292, uc_1293, uc_1294, 
      uc_1295}), .Cin(), .S({\temp1[13] [32], \temp1[13] [31], \temp1[13] [30], 
      \temp1[13] [29], \temp1[13] [28], \temp1[13] [27], \temp1[13] [26], 
      \temp1[13] [25], \temp1[13] [24], \temp1[13] [23], \temp1[13] [22], 
      \temp1[13] [21], \temp1[13] [20], \temp1[13] [19], \temp1[13] [18], 
      \temp1[13] [17], uc_1296, uc_1297, uc_1298, uc_1299, uc_1300, uc_1301, 
      uc_1302, uc_1303, uc_1304, uc_1305, uc_1306, uc_1307, uc_1308, uc_1309, 
      uc_1310, uc_1311, uc_1312}), .overFlow());
   Carry_Look_Ahead_generic__0_4908 x_13_Ux (.A({n_0_29, uc_1313, n_0_28, n_0_27, 
      n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, uc_1314, uc_1315, uc_1316, uc_1317, uc_1318, 
      uc_1319, uc_1320, uc_1321, uc_1322, uc_1323, uc_1324, uc_1325, uc_1326, 
      uc_1327, uc_1328, uc_1329, uc_1330}), .B({mn[15], mn[14], mn[13], mn[12], 
      mn[11], mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], 
      mn[1], m[0], uc_1331, uc_1332, uc_1333, uc_1334, uc_1335, uc_1336, uc_1337, 
      uc_1338, uc_1339, uc_1340, uc_1341, uc_1342, uc_1343, uc_1344, uc_1345, 
      uc_1346, uc_1347}), .Cin(), .S({\temp2[13] [32], \temp2[13] [31], 
      \temp2[13] [30], \temp2[13] [29], \temp2[13] [28], \temp2[13] [27], 
      \temp2[13] [26], \temp2[13] [25], \temp2[13] [24], \temp2[13] [23], 
      \temp2[13] [22], \temp2[13] [21], \temp2[13] [20], \temp2[13] [19], 
      \temp2[13] [18], \temp2[13] [17], uc_1348, uc_1349, uc_1350, uc_1351, 
      uc_1352, uc_1353, uc_1354, uc_1355, uc_1356, uc_1357, uc_1358, uc_1359, 
      uc_1360, uc_1361, uc_1362, uc_1363, uc_1364}), .overFlow());
   Carry_Look_Ahead_generic__0_5076 x_14_Ux (.A({n_0_14, uc_1365, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1, n_0_0, uc_1366, uc_1367, uc_1368, uc_1369, uc_1370, uc_1371, 
      uc_1372, uc_1373, uc_1374, uc_1375, uc_1376, uc_1377, uc_1378, uc_1379, 
      uc_1380, uc_1381, uc_1382}), .B({mn[15], mn[14], mn[13], mn[12], mn[11], 
      mn[10], mn[9], mn[8], mn[7], mn[6], mn[5], mn[4], mn[3], mn[2], mn[1], 
      m[0], uc_1383, uc_1384, uc_1385, uc_1386, uc_1387, uc_1388, uc_1389, 
      uc_1390, uc_1391, uc_1392, uc_1393, uc_1394, uc_1395, uc_1396, uc_1397, 
      uc_1398, uc_1399}), .Cin(), .S({\temp2[14] [32], \temp2[14] [31], 
      \temp2[14] [30], \temp2[14] [29], \temp2[14] [28], \temp2[14] [27], 
      \temp2[14] [26], \temp2[14] [25], \temp2[14] [24], \temp2[14] [23], 
      \temp2[14] [22], \temp2[14] [21], \temp2[14] [20], \temp2[14] [19], 
      \temp2[14] [18], \temp2[14] [17], uc_1400, uc_1401, uc_1402, uc_1403, 
      uc_1404, uc_1405, uc_1406, uc_1407, uc_1408, uc_1409, uc_1410, uc_1411, 
      uc_1412, uc_1413, uc_1414, uc_1415, uc_1416}), .overFlow());
   Carry_Look_Ahead_generic x_14_Un (.A({n_0_14, uc_1417, n_0_13, n_0_12, n_0_11, 
      n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, 
      n_0_0, uc_1418, uc_1419, uc_1420, uc_1421, uc_1422, uc_1423, uc_1424, 
      uc_1425, uc_1426, uc_1427, uc_1428, uc_1429, uc_1430, uc_1431, uc_1432, 
      uc_1433, uc_1434}), .B({m[15], m[14], m[13], m[12], m[11], m[10], m[9], 
      m[8], m[7], m[6], m[5], m[4], m[3], m[2], m[1], m[0], uc_1435, uc_1436, 
      uc_1437, uc_1438, uc_1439, uc_1440, uc_1441, uc_1442, uc_1443, uc_1444, 
      uc_1445, uc_1446, uc_1447, uc_1448, uc_1449, uc_1450, uc_1451}), .Cin(), 
      .S({\temp1[14] [32], \temp1[14] [31], \temp1[14] [30], \temp1[14] [29], 
      \temp1[14] [28], \temp1[14] [27], \temp1[14] [26], \temp1[14] [25], 
      \temp1[14] [24], \temp1[14] [23], \temp1[14] [22], \temp1[14] [21], 
      \temp1[14] [20], \temp1[14] [19], \temp1[14] [18], \temp1[14] [17], 
      uc_1452, uc_1453, uc_1454, uc_1455, uc_1456, uc_1457, uc_1458, uc_1459, 
      uc_1460, uc_1461, uc_1462, uc_1463, uc_1464, uc_1465, uc_1466, uc_1467, 
      uc_1468}), .overFlow());
   INV_X1 i_0_0_0 (.A(m[0]), .ZN(notM[0]));
   INV_X1 i_0_0_1 (.A(m[1]), .ZN(notM[1]));
   INV_X1 i_0_0_2 (.A(m[2]), .ZN(notM[2]));
   INV_X1 i_0_0_3 (.A(m[3]), .ZN(notM[3]));
   INV_X1 i_0_0_4 (.A(m[4]), .ZN(notM[4]));
   INV_X1 i_0_0_5 (.A(m[5]), .ZN(notM[5]));
   INV_X1 i_0_0_6 (.A(m[6]), .ZN(notM[6]));
   INV_X1 i_0_0_7 (.A(m[7]), .ZN(notM[7]));
   INV_X1 i_0_0_8 (.A(m[8]), .ZN(notM[8]));
   INV_X1 i_0_0_9 (.A(m[9]), .ZN(notM[9]));
   INV_X1 i_0_0_10 (.A(m[10]), .ZN(notM[10]));
   INV_X1 i_0_0_11 (.A(m[11]), .ZN(notM[11]));
   INV_X1 i_0_0_12 (.A(m[12]), .ZN(notM[12]));
   INV_X1 i_0_0_13 (.A(m[13]), .ZN(notM[13]));
   INV_X1 i_0_0_14 (.A(m[14]), .ZN(notM[14]));
   INV_X1 i_0_0_15 (.A(m[15]), .ZN(notM[15]));
   INV_X1 i_0_1_0 (.A(n_0_1_0), .ZN(result[0]));
   AOI222_X1 i_0_1_1 (.A1(\temp2[7] [17]), .A2(n_0_1_240), .B1(\temp1[7] [17]), 
      .B2(n_0_1_241), .C1(n_0_1_239), .C2(n_0_105), .ZN(n_0_1_0));
   INV_X1 i_0_1_2 (.A(n_0_1_1), .ZN(result[1]));
   AOI222_X1 i_0_1_3 (.A1(\temp1[8] [17]), .A2(n_0_1_235), .B1(\temp2[8] [17]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_90), .ZN(n_0_1_1));
   INV_X1 i_0_1_4 (.A(n_0_1_2), .ZN(result[2]));
   AOI222_X1 i_0_1_5 (.A1(\temp1[9] [17]), .A2(n_0_1_230), .B1(\temp2[9] [17]), 
      .B2(n_0_1_231), .C1(n_0_1_229), .C2(n_0_75), .ZN(n_0_1_2));
   INV_X1 i_0_1_6 (.A(n_0_1_3), .ZN(result[3]));
   AOI222_X1 i_0_1_7 (.A1(\temp1[10] [17]), .A2(n_0_1_225), .B1(\temp2[10] [17]), 
      .B2(n_0_1_226), .C1(n_0_1_224), .C2(n_0_60), .ZN(n_0_1_3));
   INV_X1 i_0_1_8 (.A(n_0_1_4), .ZN(result[4]));
   AOI222_X1 i_0_1_9 (.A1(\temp1[11] [17]), .A2(n_0_1_220), .B1(\temp2[11] [17]), 
      .B2(n_0_1_221), .C1(n_0_1_219), .C2(n_0_45), .ZN(n_0_1_4));
   INV_X1 i_0_1_10 (.A(n_0_1_5), .ZN(result[5]));
   AOI222_X1 i_0_1_11 (.A1(\temp1[12] [17]), .A2(n_0_1_216), .B1(\temp2[12] [17]), 
      .B2(n_0_1_215), .C1(n_0_1_214), .C2(n_0_30), .ZN(n_0_1_5));
   INV_X1 i_0_1_12 (.A(n_0_1_6), .ZN(result[6]));
   AOI222_X1 i_0_1_13 (.A1(\temp2[13] [17]), .A2(n_0_1_274), .B1(\temp1[13] [17]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_15), .ZN(n_0_1_6));
   INV_X1 i_0_1_14 (.A(n_0_1_7), .ZN(result[7]));
   AOI222_X1 i_0_1_15 (.A1(\temp1[14] [17]), .A2(n_0_1_277), .B1(\temp2[14] [17]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_0), .ZN(n_0_1_7));
   INV_X1 i_0_1_16 (.A(n_0_1_8), .ZN(result[8]));
   AOI222_X1 i_0_1_17 (.A1(\temp1[14] [18]), .A2(n_0_1_277), .B1(\temp2[14] [18]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_1), .ZN(n_0_1_8));
   INV_X1 i_0_1_18 (.A(n_0_1_9), .ZN(result[9]));
   AOI222_X1 i_0_1_19 (.A1(\temp1[14] [19]), .A2(n_0_1_277), .B1(\temp2[14] [19]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_2), .ZN(n_0_1_9));
   INV_X1 i_0_1_20 (.A(n_0_1_10), .ZN(result[10]));
   AOI222_X1 i_0_1_21 (.A1(\temp1[14] [20]), .A2(n_0_1_277), .B1(\temp2[14] [20]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_3), .ZN(n_0_1_10));
   INV_X1 i_0_1_22 (.A(n_0_1_11), .ZN(result[11]));
   AOI222_X1 i_0_1_23 (.A1(\temp1[14] [21]), .A2(n_0_1_277), .B1(\temp2[14] [21]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_4), .ZN(n_0_1_11));
   INV_X1 i_0_1_24 (.A(n_0_1_12), .ZN(result[12]));
   AOI222_X1 i_0_1_25 (.A1(\temp1[14] [22]), .A2(n_0_1_277), .B1(\temp2[14] [22]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_5), .ZN(n_0_1_12));
   INV_X1 i_0_1_26 (.A(n_0_1_13), .ZN(result[13]));
   AOI222_X1 i_0_1_27 (.A1(\temp1[14] [23]), .A2(n_0_1_277), .B1(\temp2[14] [23]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_6), .ZN(n_0_1_13));
   INV_X1 i_0_1_28 (.A(n_0_1_14), .ZN(result[14]));
   AOI222_X1 i_0_1_29 (.A1(\temp1[14] [24]), .A2(n_0_1_277), .B1(\temp2[14] [24]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_7), .ZN(n_0_1_14));
   INV_X1 i_0_1_30 (.A(n_0_1_15), .ZN(result[15]));
   AOI222_X1 i_0_1_31 (.A1(\temp1[14] [25]), .A2(n_0_1_277), .B1(\temp2[14] [25]), 
      .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_8), .ZN(n_0_1_15));
   INV_X1 i_0_1_32 (.A(n_0_1_16), .ZN(n_0_0));
   AOI222_X1 i_0_1_33 (.A1(\temp2[13] [18]), .A2(n_0_1_274), .B1(\temp1[13] [18]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_16), .ZN(n_0_1_16));
   INV_X1 i_0_1_34 (.A(n_0_1_17), .ZN(n_0_1));
   AOI222_X1 i_0_1_35 (.A1(\temp2[13] [19]), .A2(n_0_1_274), .B1(\temp1[13] [19]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_17), .ZN(n_0_1_17));
   INV_X1 i_0_1_36 (.A(n_0_1_18), .ZN(n_0_2));
   AOI222_X1 i_0_1_37 (.A1(\temp2[13] [20]), .A2(n_0_1_274), .B1(\temp1[13] [20]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_18), .ZN(n_0_1_18));
   INV_X1 i_0_1_38 (.A(n_0_1_19), .ZN(n_0_3));
   AOI222_X1 i_0_1_39 (.A1(\temp2[13] [21]), .A2(n_0_1_274), .B1(\temp1[13] [21]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_19), .ZN(n_0_1_19));
   INV_X1 i_0_1_40 (.A(n_0_1_20), .ZN(n_0_4));
   AOI222_X1 i_0_1_41 (.A1(\temp2[13] [22]), .A2(n_0_1_274), .B1(\temp1[13] [22]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_20), .ZN(n_0_1_20));
   INV_X1 i_0_1_42 (.A(n_0_1_21), .ZN(n_0_5));
   AOI222_X1 i_0_1_43 (.A1(\temp2[13] [23]), .A2(n_0_1_274), .B1(\temp1[13] [23]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_21), .ZN(n_0_1_21));
   INV_X1 i_0_1_44 (.A(n_0_1_22), .ZN(n_0_6));
   AOI222_X1 i_0_1_45 (.A1(\temp2[13] [24]), .A2(n_0_1_274), .B1(\temp1[13] [24]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_22), .ZN(n_0_1_22));
   INV_X1 i_0_1_46 (.A(n_0_1_23), .ZN(n_0_7));
   AOI222_X1 i_0_1_47 (.A1(\temp2[13] [25]), .A2(n_0_1_274), .B1(\temp1[13] [25]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_23), .ZN(n_0_1_23));
   INV_X1 i_0_1_48 (.A(n_0_1_24), .ZN(n_0_8));
   AOI222_X1 i_0_1_49 (.A1(\temp2[13] [26]), .A2(n_0_1_274), .B1(\temp1[13] [26]), 
      .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_24), .ZN(n_0_1_24));
   INV_X1 i_0_1_50 (.A(n_0_1_25), .ZN(n_0_15));
   AOI222_X1 i_0_1_51 (.A1(\temp1[12] [18]), .A2(n_0_1_216), .B1(\temp2[12] [18]), 
      .B2(n_0_1_215), .C1(n_0_1_214), .C2(n_0_31), .ZN(n_0_1_25));
   INV_X1 i_0_1_52 (.A(n_0_1_26), .ZN(n_0_16));
   AOI222_X1 i_0_1_53 (.A1(\temp2[12] [19]), .A2(n_0_1_215), .B1(\temp1[12] [19]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_32), .ZN(n_0_1_26));
   INV_X1 i_0_1_54 (.A(n_0_1_27), .ZN(n_0_17));
   AOI222_X1 i_0_1_55 (.A1(\temp2[12] [20]), .A2(n_0_1_215), .B1(\temp1[12] [20]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_33), .ZN(n_0_1_27));
   INV_X1 i_0_1_56 (.A(n_0_1_28), .ZN(n_0_18));
   AOI222_X1 i_0_1_57 (.A1(\temp2[12] [21]), .A2(n_0_1_215), .B1(\temp1[12] [21]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_34), .ZN(n_0_1_28));
   INV_X1 i_0_1_58 (.A(n_0_1_29), .ZN(n_0_19));
   AOI222_X1 i_0_1_59 (.A1(\temp2[12] [22]), .A2(n_0_1_215), .B1(\temp1[12] [22]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_35), .ZN(n_0_1_29));
   INV_X1 i_0_1_60 (.A(n_0_1_30), .ZN(n_0_20));
   AOI222_X1 i_0_1_61 (.A1(\temp2[12] [23]), .A2(n_0_1_215), .B1(\temp1[12] [23]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_36), .ZN(n_0_1_30));
   INV_X1 i_0_1_62 (.A(n_0_1_31), .ZN(n_0_21));
   AOI222_X1 i_0_1_63 (.A1(\temp2[12] [24]), .A2(n_0_1_215), .B1(\temp1[12] [24]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_37), .ZN(n_0_1_31));
   INV_X1 i_0_1_64 (.A(n_0_1_32), .ZN(n_0_22));
   AOI222_X1 i_0_1_65 (.A1(\temp2[12] [25]), .A2(n_0_1_215), .B1(\temp1[12] [25]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_38), .ZN(n_0_1_32));
   INV_X1 i_0_1_66 (.A(n_0_1_33), .ZN(n_0_23));
   AOI222_X1 i_0_1_67 (.A1(\temp2[12] [26]), .A2(n_0_1_215), .B1(\temp1[12] [26]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_39), .ZN(n_0_1_33));
   INV_X1 i_0_1_68 (.A(n_0_1_34), .ZN(n_0_24));
   AOI222_X1 i_0_1_69 (.A1(\temp2[12] [27]), .A2(n_0_1_215), .B1(\temp1[12] [27]), 
      .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_40), .ZN(n_0_1_34));
   INV_X1 i_0_1_70 (.A(n_0_1_35), .ZN(n_0_30));
   AOI222_X1 i_0_1_71 (.A1(\temp2[11] [18]), .A2(n_0_1_221), .B1(\temp1[11] [18]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_46), .ZN(n_0_1_35));
   INV_X1 i_0_1_72 (.A(n_0_1_36), .ZN(n_0_31));
   AOI222_X1 i_0_1_73 (.A1(\temp2[11] [19]), .A2(n_0_1_221), .B1(\temp1[11] [19]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_47), .ZN(n_0_1_36));
   INV_X1 i_0_1_74 (.A(n_0_1_37), .ZN(n_0_32));
   AOI222_X1 i_0_1_75 (.A1(\temp2[11] [20]), .A2(n_0_1_221), .B1(\temp1[11] [20]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_48), .ZN(n_0_1_37));
   INV_X1 i_0_1_76 (.A(n_0_1_38), .ZN(n_0_33));
   AOI222_X1 i_0_1_77 (.A1(\temp2[11] [21]), .A2(n_0_1_221), .B1(\temp1[11] [21]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_49), .ZN(n_0_1_38));
   INV_X1 i_0_1_78 (.A(n_0_1_39), .ZN(n_0_34));
   AOI222_X1 i_0_1_79 (.A1(\temp2[11] [22]), .A2(n_0_1_221), .B1(\temp1[11] [22]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_50), .ZN(n_0_1_39));
   INV_X1 i_0_1_80 (.A(n_0_1_40), .ZN(n_0_35));
   AOI222_X1 i_0_1_81 (.A1(\temp2[11] [23]), .A2(n_0_1_221), .B1(\temp1[11] [23]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_51), .ZN(n_0_1_40));
   INV_X1 i_0_1_82 (.A(n_0_1_41), .ZN(n_0_36));
   AOI222_X1 i_0_1_83 (.A1(\temp2[11] [24]), .A2(n_0_1_221), .B1(\temp1[11] [24]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_52), .ZN(n_0_1_41));
   INV_X1 i_0_1_84 (.A(n_0_1_42), .ZN(n_0_37));
   AOI222_X1 i_0_1_85 (.A1(\temp2[11] [25]), .A2(n_0_1_221), .B1(\temp1[11] [25]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_53), .ZN(n_0_1_42));
   INV_X1 i_0_1_86 (.A(n_0_1_43), .ZN(n_0_38));
   AOI222_X1 i_0_1_87 (.A1(\temp2[11] [26]), .A2(n_0_1_221), .B1(\temp1[11] [26]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_54), .ZN(n_0_1_43));
   INV_X1 i_0_1_88 (.A(n_0_1_44), .ZN(n_0_39));
   AOI222_X1 i_0_1_89 (.A1(\temp2[11] [27]), .A2(n_0_1_221), .B1(\temp1[11] [27]), 
      .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_55), .ZN(n_0_1_44));
   INV_X1 i_0_1_90 (.A(n_0_1_45), .ZN(n_0_40));
   AOI222_X1 i_0_1_91 (.A1(\temp1[11] [28]), .A2(n_0_1_220), .B1(\temp2[11] [28]), 
      .B2(n_0_1_221), .C1(n_0_1_219), .C2(n_0_56), .ZN(n_0_1_45));
   INV_X1 i_0_1_92 (.A(n_0_1_46), .ZN(n_0_45));
   AOI222_X1 i_0_1_93 (.A1(\temp1[10] [18]), .A2(n_0_1_225), .B1(\temp2[10] [18]), 
      .B2(n_0_1_226), .C1(n_0_1_224), .C2(n_0_61), .ZN(n_0_1_46));
   INV_X1 i_0_1_94 (.A(n_0_1_47), .ZN(n_0_46));
   AOI222_X1 i_0_1_95 (.A1(\temp2[10] [19]), .A2(n_0_1_226), .B1(\temp1[10] [19]), 
      .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_62), .ZN(n_0_1_47));
   INV_X1 i_0_1_96 (.A(n_0_1_48), .ZN(n_0_47));
   AOI222_X1 i_0_1_97 (.A1(\temp2[10] [20]), .A2(n_0_1_226), .B1(\temp1[10] [20]), 
      .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_63), .ZN(n_0_1_48));
   INV_X1 i_0_1_98 (.A(n_0_1_49), .ZN(n_0_48));
   AOI222_X1 i_0_1_99 (.A1(\temp2[10] [21]), .A2(n_0_1_226), .B1(\temp1[10] [21]), 
      .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_64), .ZN(n_0_1_49));
   INV_X1 i_0_1_100 (.A(n_0_1_50), .ZN(n_0_49));
   AOI222_X1 i_0_1_101 (.A1(\temp2[10] [22]), .A2(n_0_1_226), .B1(
      \temp1[10] [22]), .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_65), .ZN(
      n_0_1_50));
   INV_X1 i_0_1_102 (.A(n_0_1_51), .ZN(n_0_50));
   AOI222_X1 i_0_1_103 (.A1(\temp2[10] [23]), .A2(n_0_1_226), .B1(
      \temp1[10] [23]), .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_66), .ZN(
      n_0_1_51));
   INV_X1 i_0_1_104 (.A(n_0_1_52), .ZN(n_0_51));
   AOI222_X1 i_0_1_105 (.A1(\temp2[10] [24]), .A2(n_0_1_226), .B1(
      \temp1[10] [24]), .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_67), .ZN(
      n_0_1_52));
   INV_X1 i_0_1_106 (.A(n_0_1_53), .ZN(n_0_52));
   AOI222_X1 i_0_1_107 (.A1(\temp2[10] [25]), .A2(n_0_1_226), .B1(
      \temp1[10] [25]), .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_68), .ZN(
      n_0_1_53));
   INV_X1 i_0_1_108 (.A(n_0_1_54), .ZN(n_0_53));
   AOI222_X1 i_0_1_109 (.A1(\temp2[10] [26]), .A2(n_0_1_226), .B1(
      \temp1[10] [26]), .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_69), .ZN(
      n_0_1_54));
   INV_X1 i_0_1_110 (.A(n_0_1_55), .ZN(n_0_54));
   AOI222_X1 i_0_1_111 (.A1(\temp2[10] [27]), .A2(n_0_1_226), .B1(
      \temp1[10] [27]), .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_70), .ZN(
      n_0_1_55));
   INV_X1 i_0_1_112 (.A(n_0_1_56), .ZN(n_0_55));
   AOI222_X1 i_0_1_113 (.A1(\temp1[10] [28]), .A2(n_0_1_225), .B1(
      \temp2[10] [28]), .B2(n_0_1_226), .C1(n_0_1_224), .C2(n_0_71), .ZN(
      n_0_1_56));
   INV_X1 i_0_1_114 (.A(n_0_1_57), .ZN(n_0_56));
   AOI222_X1 i_0_1_115 (.A1(\temp1[10] [29]), .A2(n_0_1_225), .B1(
      \temp2[10] [29]), .B2(n_0_1_226), .C1(n_0_1_224), .C2(n_0_72), .ZN(
      n_0_1_57));
   INV_X1 i_0_1_116 (.A(n_0_1_58), .ZN(n_0_60));
   AOI222_X1 i_0_1_117 (.A1(\temp1[9] [18]), .A2(n_0_1_230), .B1(\temp2[9] [18]), 
      .B2(n_0_1_231), .C1(n_0_1_229), .C2(n_0_76), .ZN(n_0_1_58));
   INV_X1 i_0_1_118 (.A(n_0_1_59), .ZN(n_0_61));
   AOI222_X1 i_0_1_119 (.A1(\temp1[9] [19]), .A2(n_0_1_230), .B1(\temp2[9] [19]), 
      .B2(n_0_1_231), .C1(n_0_1_229), .C2(n_0_77), .ZN(n_0_1_59));
   INV_X1 i_0_1_120 (.A(n_0_1_60), .ZN(n_0_62));
   AOI222_X1 i_0_1_121 (.A1(\temp1[9] [20]), .A2(n_0_1_230), .B1(\temp2[9] [20]), 
      .B2(n_0_1_231), .C1(n_0_1_229), .C2(n_0_78), .ZN(n_0_1_60));
   INV_X1 i_0_1_122 (.A(n_0_1_61), .ZN(n_0_63));
   AOI222_X1 i_0_1_123 (.A1(\temp2[9] [21]), .A2(n_0_1_231), .B1(\temp1[9] [21]), 
      .B2(n_0_1_230), .C1(n_0_1_229), .C2(n_0_79), .ZN(n_0_1_61));
   INV_X1 i_0_1_124 (.A(n_0_1_62), .ZN(n_0_64));
   AOI222_X1 i_0_1_125 (.A1(\temp2[9] [22]), .A2(n_0_1_231), .B1(\temp1[9] [22]), 
      .B2(n_0_1_230), .C1(n_0_1_229), .C2(n_0_80), .ZN(n_0_1_62));
   INV_X1 i_0_1_126 (.A(n_0_1_63), .ZN(n_0_65));
   AOI222_X1 i_0_1_127 (.A1(\temp2[9] [23]), .A2(n_0_1_231), .B1(\temp1[9] [23]), 
      .B2(n_0_1_230), .C1(n_0_1_229), .C2(n_0_81), .ZN(n_0_1_63));
   INV_X1 i_0_1_128 (.A(n_0_1_64), .ZN(n_0_66));
   AOI222_X1 i_0_1_129 (.A1(\temp2[9] [24]), .A2(n_0_1_231), .B1(\temp1[9] [24]), 
      .B2(n_0_1_230), .C1(n_0_1_229), .C2(n_0_82), .ZN(n_0_1_64));
   INV_X1 i_0_1_130 (.A(n_0_1_65), .ZN(n_0_67));
   AOI222_X1 i_0_1_131 (.A1(\temp2[9] [25]), .A2(n_0_1_231), .B1(\temp1[9] [25]), 
      .B2(n_0_1_230), .C1(n_0_1_229), .C2(n_0_83), .ZN(n_0_1_65));
   INV_X1 i_0_1_132 (.A(n_0_1_66), .ZN(n_0_68));
   AOI222_X1 i_0_1_133 (.A1(\temp2[9] [26]), .A2(n_0_1_231), .B1(\temp1[9] [26]), 
      .B2(n_0_1_230), .C1(n_0_1_229), .C2(n_0_84), .ZN(n_0_1_66));
   INV_X1 i_0_1_134 (.A(n_0_1_67), .ZN(n_0_69));
   AOI222_X1 i_0_1_135 (.A1(\temp2[9] [27]), .A2(n_0_1_231), .B1(\temp1[9] [27]), 
      .B2(n_0_1_230), .C1(n_0_1_229), .C2(n_0_85), .ZN(n_0_1_67));
   INV_X1 i_0_1_136 (.A(n_0_1_68), .ZN(n_0_70));
   AOI222_X1 i_0_1_137 (.A1(\temp1[9] [28]), .A2(n_0_1_230), .B1(\temp2[9] [28]), 
      .B2(n_0_1_231), .C1(n_0_1_229), .C2(n_0_86), .ZN(n_0_1_68));
   INV_X1 i_0_1_138 (.A(n_0_1_69), .ZN(n_0_71));
   AOI222_X1 i_0_1_139 (.A1(\temp1[9] [29]), .A2(n_0_1_230), .B1(\temp2[9] [29]), 
      .B2(n_0_1_231), .C1(n_0_1_229), .C2(n_0_87), .ZN(n_0_1_69));
   INV_X1 i_0_1_140 (.A(n_0_1_70), .ZN(n_0_72));
   AOI222_X1 i_0_1_141 (.A1(\temp1[9] [30]), .A2(n_0_1_230), .B1(\temp2[9] [30]), 
      .B2(n_0_1_231), .C1(n_0_1_229), .C2(n_0_88), .ZN(n_0_1_70));
   INV_X1 i_0_1_142 (.A(n_0_1_71), .ZN(n_0_75));
   AOI222_X1 i_0_1_143 (.A1(\temp1[8] [18]), .A2(n_0_1_235), .B1(\temp2[8] [18]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_91), .ZN(n_0_1_71));
   INV_X1 i_0_1_144 (.A(n_0_1_72), .ZN(n_0_76));
   AOI222_X1 i_0_1_145 (.A1(\temp1[8] [19]), .A2(n_0_1_235), .B1(\temp2[8] [19]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_92), .ZN(n_0_1_72));
   INV_X1 i_0_1_146 (.A(n_0_1_73), .ZN(n_0_77));
   AOI222_X1 i_0_1_147 (.A1(\temp1[8] [20]), .A2(n_0_1_235), .B1(\temp2[8] [20]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_93), .ZN(n_0_1_73));
   INV_X1 i_0_1_148 (.A(n_0_1_74), .ZN(n_0_78));
   AOI222_X1 i_0_1_149 (.A1(\temp1[8] [21]), .A2(n_0_1_235), .B1(\temp2[8] [21]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_94), .ZN(n_0_1_74));
   INV_X1 i_0_1_150 (.A(n_0_1_75), .ZN(n_0_79));
   AOI222_X1 i_0_1_151 (.A1(\temp2[8] [22]), .A2(n_0_1_236), .B1(\temp1[8] [22]), 
      .B2(n_0_1_235), .C1(n_0_1_234), .C2(n_0_95), .ZN(n_0_1_75));
   INV_X1 i_0_1_152 (.A(n_0_1_76), .ZN(n_0_80));
   AOI222_X1 i_0_1_153 (.A1(\temp2[8] [23]), .A2(n_0_1_236), .B1(\temp1[8] [23]), 
      .B2(n_0_1_235), .C1(n_0_1_234), .C2(n_0_96), .ZN(n_0_1_76));
   INV_X1 i_0_1_154 (.A(n_0_1_77), .ZN(n_0_81));
   AOI222_X1 i_0_1_155 (.A1(\temp2[8] [24]), .A2(n_0_1_236), .B1(\temp1[8] [24]), 
      .B2(n_0_1_235), .C1(n_0_1_234), .C2(n_0_97), .ZN(n_0_1_77));
   INV_X1 i_0_1_156 (.A(n_0_1_78), .ZN(n_0_82));
   AOI222_X1 i_0_1_157 (.A1(\temp2[8] [25]), .A2(n_0_1_236), .B1(\temp1[8] [25]), 
      .B2(n_0_1_235), .C1(n_0_1_234), .C2(n_0_98), .ZN(n_0_1_78));
   INV_X1 i_0_1_158 (.A(n_0_1_79), .ZN(n_0_83));
   AOI222_X1 i_0_1_159 (.A1(\temp2[8] [26]), .A2(n_0_1_236), .B1(\temp1[8] [26]), 
      .B2(n_0_1_235), .C1(n_0_1_234), .C2(n_0_99), .ZN(n_0_1_79));
   INV_X1 i_0_1_160 (.A(n_0_1_80), .ZN(n_0_84));
   AOI222_X1 i_0_1_161 (.A1(\temp2[8] [27]), .A2(n_0_1_236), .B1(\temp1[8] [27]), 
      .B2(n_0_1_235), .C1(n_0_1_234), .C2(n_0_100), .ZN(n_0_1_80));
   INV_X1 i_0_1_162 (.A(n_0_1_81), .ZN(n_0_85));
   AOI222_X1 i_0_1_163 (.A1(\temp1[8] [28]), .A2(n_0_1_235), .B1(\temp2[8] [28]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_101), .ZN(n_0_1_81));
   INV_X1 i_0_1_164 (.A(n_0_1_82), .ZN(n_0_86));
   AOI222_X1 i_0_1_165 (.A1(\temp1[8] [29]), .A2(n_0_1_235), .B1(\temp2[8] [29]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_102), .ZN(n_0_1_82));
   INV_X1 i_0_1_166 (.A(n_0_1_83), .ZN(n_0_87));
   AOI222_X1 i_0_1_167 (.A1(\temp1[8] [30]), .A2(n_0_1_235), .B1(\temp2[8] [30]), 
      .B2(n_0_1_236), .C1(n_0_1_234), .C2(n_0_103), .ZN(n_0_1_83));
   INV_X1 i_0_1_168 (.A(n_0_1_84), .ZN(n_0_88));
   AOI221_X1 i_0_1_169 (.A(n_0_1_233), .B1(\temp2[8] [31]), .B2(n_0_1_236), 
      .C1(\temp1[8] [31]), .C2(n_0_1_235), .ZN(n_0_1_84));
   INV_X1 i_0_1_170 (.A(n_0_1_85), .ZN(n_0_90));
   AOI222_X1 i_0_1_171 (.A1(\temp2[7] [18]), .A2(n_0_1_240), .B1(\temp1[7] [18]), 
      .B2(n_0_1_241), .C1(n_0_1_239), .C2(n_0_106), .ZN(n_0_1_85));
   INV_X1 i_0_1_172 (.A(n_0_1_86), .ZN(n_0_91));
   AOI222_X1 i_0_1_173 (.A1(\temp1[7] [19]), .A2(n_0_1_241), .B1(\temp2[7] [19]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_107), .ZN(n_0_1_86));
   INV_X1 i_0_1_174 (.A(n_0_1_87), .ZN(n_0_92));
   AOI222_X1 i_0_1_175 (.A1(\temp1[7] [20]), .A2(n_0_1_241), .B1(\temp2[7] [20]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_108), .ZN(n_0_1_87));
   INV_X1 i_0_1_176 (.A(n_0_1_88), .ZN(n_0_93));
   AOI222_X1 i_0_1_177 (.A1(\temp1[7] [21]), .A2(n_0_1_241), .B1(\temp2[7] [21]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_109), .ZN(n_0_1_88));
   INV_X1 i_0_1_178 (.A(n_0_1_89), .ZN(n_0_94));
   AOI222_X1 i_0_1_179 (.A1(\temp1[7] [22]), .A2(n_0_1_241), .B1(\temp2[7] [22]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_110), .ZN(n_0_1_89));
   INV_X1 i_0_1_180 (.A(n_0_1_90), .ZN(n_0_95));
   AOI222_X1 i_0_1_181 (.A1(\temp1[7] [23]), .A2(n_0_1_241), .B1(\temp2[7] [23]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_111), .ZN(n_0_1_90));
   INV_X1 i_0_1_182 (.A(n_0_1_91), .ZN(n_0_96));
   AOI222_X1 i_0_1_183 (.A1(\temp2[7] [24]), .A2(n_0_1_240), .B1(\temp1[7] [24]), 
      .B2(n_0_1_241), .C1(n_0_1_239), .C2(n_0_112), .ZN(n_0_1_91));
   INV_X1 i_0_1_184 (.A(n_0_1_92), .ZN(n_0_97));
   AOI222_X1 i_0_1_185 (.A1(\temp2[7] [25]), .A2(n_0_1_240), .B1(\temp1[7] [25]), 
      .B2(n_0_1_241), .C1(n_0_1_239), .C2(n_0_113), .ZN(n_0_1_92));
   INV_X1 i_0_1_186 (.A(n_0_1_93), .ZN(n_0_98));
   AOI222_X1 i_0_1_187 (.A1(\temp2[7] [26]), .A2(n_0_1_240), .B1(\temp1[7] [26]), 
      .B2(n_0_1_241), .C1(n_0_1_239), .C2(n_0_114), .ZN(n_0_1_93));
   INV_X1 i_0_1_188 (.A(n_0_1_94), .ZN(n_0_99));
   AOI222_X1 i_0_1_189 (.A1(\temp2[7] [27]), .A2(n_0_1_240), .B1(\temp1[7] [27]), 
      .B2(n_0_1_241), .C1(n_0_1_239), .C2(n_0_115), .ZN(n_0_1_94));
   INV_X1 i_0_1_190 (.A(n_0_1_95), .ZN(n_0_100));
   AOI222_X1 i_0_1_191 (.A1(\temp1[7] [28]), .A2(n_0_1_241), .B1(\temp2[7] [28]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_116), .ZN(n_0_1_95));
   INV_X1 i_0_1_192 (.A(n_0_1_96), .ZN(n_0_101));
   AOI222_X1 i_0_1_193 (.A1(\temp1[7] [29]), .A2(n_0_1_241), .B1(\temp2[7] [29]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_117), .ZN(n_0_1_96));
   INV_X1 i_0_1_194 (.A(n_0_1_97), .ZN(n_0_102));
   AOI222_X1 i_0_1_195 (.A1(\temp1[7] [30]), .A2(n_0_1_241), .B1(\temp2[7] [30]), 
      .B2(n_0_1_240), .C1(n_0_1_239), .C2(n_0_118), .ZN(n_0_1_97));
   INV_X1 i_0_1_196 (.A(n_0_1_98), .ZN(n_0_103));
   AOI221_X1 i_0_1_197 (.A(n_0_1_238), .B1(\temp2[7] [31]), .B2(n_0_1_240), 
      .C1(\temp1[7] [31]), .C2(n_0_1_241), .ZN(n_0_1_98));
   INV_X1 i_0_1_198 (.A(n_0_1_99), .ZN(n_0_105));
   AOI222_X1 i_0_1_199 (.A1(\temp1[6] [18]), .A2(n_0_1_245), .B1(\temp2[6] [18]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_121), .ZN(n_0_1_99));
   INV_X1 i_0_1_200 (.A(n_0_1_100), .ZN(n_0_106));
   AOI222_X1 i_0_1_201 (.A1(\temp1[6] [19]), .A2(n_0_1_245), .B1(\temp2[6] [19]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_122), .ZN(n_0_1_100));
   INV_X1 i_0_1_202 (.A(n_0_1_101), .ZN(n_0_107));
   AOI222_X1 i_0_1_203 (.A1(\temp1[6] [20]), .A2(n_0_1_245), .B1(\temp2[6] [20]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_123), .ZN(n_0_1_101));
   INV_X1 i_0_1_204 (.A(n_0_1_102), .ZN(n_0_108));
   AOI222_X1 i_0_1_205 (.A1(\temp1[6] [21]), .A2(n_0_1_245), .B1(\temp2[6] [21]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_124), .ZN(n_0_1_102));
   INV_X1 i_0_1_206 (.A(n_0_1_103), .ZN(n_0_109));
   AOI222_X1 i_0_1_207 (.A1(\temp1[6] [22]), .A2(n_0_1_245), .B1(\temp2[6] [22]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_125), .ZN(n_0_1_103));
   INV_X1 i_0_1_208 (.A(n_0_1_104), .ZN(n_0_110));
   AOI222_X1 i_0_1_209 (.A1(\temp1[6] [23]), .A2(n_0_1_245), .B1(\temp2[6] [23]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_126), .ZN(n_0_1_104));
   INV_X1 i_0_1_210 (.A(n_0_1_105), .ZN(n_0_111));
   AOI222_X1 i_0_1_211 (.A1(\temp1[6] [24]), .A2(n_0_1_245), .B1(\temp2[6] [24]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_127), .ZN(n_0_1_105));
   INV_X1 i_0_1_212 (.A(n_0_1_106), .ZN(n_0_112));
   AOI222_X1 i_0_1_213 (.A1(\temp2[6] [25]), .A2(n_0_1_246), .B1(\temp1[6] [25]), 
      .B2(n_0_1_245), .C1(n_0_1_244), .C2(n_0_128), .ZN(n_0_1_106));
   INV_X1 i_0_1_214 (.A(n_0_1_107), .ZN(n_0_113));
   AOI222_X1 i_0_1_215 (.A1(\temp2[6] [26]), .A2(n_0_1_246), .B1(\temp1[6] [26]), 
      .B2(n_0_1_245), .C1(n_0_1_244), .C2(n_0_129), .ZN(n_0_1_107));
   INV_X1 i_0_1_216 (.A(n_0_1_108), .ZN(n_0_114));
   AOI222_X1 i_0_1_217 (.A1(\temp2[6] [27]), .A2(n_0_1_246), .B1(\temp1[6] [27]), 
      .B2(n_0_1_245), .C1(n_0_1_244), .C2(n_0_130), .ZN(n_0_1_108));
   INV_X1 i_0_1_218 (.A(n_0_1_109), .ZN(n_0_115));
   AOI222_X1 i_0_1_219 (.A1(\temp1[6] [28]), .A2(n_0_1_245), .B1(\temp2[6] [28]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_131), .ZN(n_0_1_109));
   INV_X1 i_0_1_220 (.A(n_0_1_110), .ZN(n_0_116));
   AOI222_X1 i_0_1_221 (.A1(\temp1[6] [29]), .A2(n_0_1_245), .B1(\temp2[6] [29]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_132), .ZN(n_0_1_110));
   INV_X1 i_0_1_222 (.A(n_0_1_111), .ZN(n_0_117));
   AOI222_X1 i_0_1_223 (.A1(\temp1[6] [30]), .A2(n_0_1_245), .B1(\temp2[6] [30]), 
      .B2(n_0_1_246), .C1(n_0_1_244), .C2(n_0_133), .ZN(n_0_1_111));
   INV_X1 i_0_1_224 (.A(n_0_1_112), .ZN(n_0_118));
   AOI221_X1 i_0_1_225 (.A(n_0_1_243), .B1(\temp2[6] [31]), .B2(n_0_1_246), 
      .C1(\temp1[6] [31]), .C2(n_0_1_245), .ZN(n_0_1_112));
   INV_X1 i_0_1_226 (.A(n_0_1_113), .ZN(n_0_120));
   AOI222_X1 i_0_1_227 (.A1(\temp1[5] [18]), .A2(n_0_1_250), .B1(\temp2[5] [18]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_136), .ZN(n_0_1_113));
   INV_X1 i_0_1_228 (.A(n_0_1_114), .ZN(n_0_121));
   AOI222_X1 i_0_1_229 (.A1(\temp1[5] [19]), .A2(n_0_1_250), .B1(\temp2[5] [19]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_137), .ZN(n_0_1_114));
   INV_X1 i_0_1_230 (.A(n_0_1_115), .ZN(n_0_122));
   AOI222_X1 i_0_1_231 (.A1(\temp1[5] [20]), .A2(n_0_1_250), .B1(\temp2[5] [20]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_138), .ZN(n_0_1_115));
   INV_X1 i_0_1_232 (.A(n_0_1_116), .ZN(n_0_123));
   AOI222_X1 i_0_1_233 (.A1(\temp1[5] [21]), .A2(n_0_1_250), .B1(\temp2[5] [21]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_139), .ZN(n_0_1_116));
   INV_X1 i_0_1_234 (.A(n_0_1_117), .ZN(n_0_124));
   AOI222_X1 i_0_1_235 (.A1(\temp1[5] [22]), .A2(n_0_1_250), .B1(\temp2[5] [22]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_140), .ZN(n_0_1_117));
   INV_X1 i_0_1_236 (.A(n_0_1_118), .ZN(n_0_125));
   AOI222_X1 i_0_1_237 (.A1(\temp1[5] [23]), .A2(n_0_1_250), .B1(\temp2[5] [23]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_141), .ZN(n_0_1_118));
   INV_X1 i_0_1_238 (.A(n_0_1_119), .ZN(n_0_126));
   AOI222_X1 i_0_1_239 (.A1(\temp1[5] [24]), .A2(n_0_1_250), .B1(\temp2[5] [24]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_142), .ZN(n_0_1_119));
   INV_X1 i_0_1_240 (.A(n_0_1_120), .ZN(n_0_127));
   AOI222_X1 i_0_1_241 (.A1(\temp1[5] [25]), .A2(n_0_1_250), .B1(\temp2[5] [25]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_143), .ZN(n_0_1_120));
   INV_X1 i_0_1_242 (.A(n_0_1_121), .ZN(n_0_128));
   AOI222_X1 i_0_1_243 (.A1(\temp1[5] [26]), .A2(n_0_1_250), .B1(\temp2[5] [26]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_144), .ZN(n_0_1_121));
   INV_X1 i_0_1_244 (.A(n_0_1_122), .ZN(n_0_129));
   AOI222_X1 i_0_1_245 (.A1(\temp1[5] [27]), .A2(n_0_1_250), .B1(\temp2[5] [27]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_145), .ZN(n_0_1_122));
   INV_X1 i_0_1_246 (.A(n_0_1_123), .ZN(n_0_130));
   AOI222_X1 i_0_1_247 (.A1(\temp1[5] [28]), .A2(n_0_1_250), .B1(\temp2[5] [28]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_146), .ZN(n_0_1_123));
   INV_X1 i_0_1_248 (.A(n_0_1_124), .ZN(n_0_131));
   AOI222_X1 i_0_1_249 (.A1(\temp1[5] [29]), .A2(n_0_1_250), .B1(\temp2[5] [29]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_147), .ZN(n_0_1_124));
   INV_X1 i_0_1_250 (.A(n_0_1_125), .ZN(n_0_132));
   AOI222_X1 i_0_1_251 (.A1(\temp1[5] [30]), .A2(n_0_1_250), .B1(\temp2[5] [30]), 
      .B2(n_0_1_251), .C1(n_0_1_249), .C2(n_0_148), .ZN(n_0_1_125));
   INV_X1 i_0_1_252 (.A(n_0_1_126), .ZN(n_0_133));
   AOI221_X1 i_0_1_253 (.A(n_0_1_248), .B1(\temp2[5] [31]), .B2(n_0_1_251), 
      .C1(\temp1[5] [31]), .C2(n_0_1_250), .ZN(n_0_1_126));
   INV_X1 i_0_1_254 (.A(n_0_1_127), .ZN(n_0_135));
   AOI222_X1 i_0_1_255 (.A1(\temp2[4] [18]), .A2(n_0_1_255), .B1(\temp1[4] [18]), 
      .B2(n_0_1_256), .C1(n_0_1_254), .C2(n_0_151), .ZN(n_0_1_127));
   INV_X1 i_0_1_256 (.A(n_0_1_128), .ZN(n_0_136));
   AOI222_X1 i_0_1_257 (.A1(\temp2[4] [19]), .A2(n_0_1_255), .B1(\temp1[4] [19]), 
      .B2(n_0_1_256), .C1(n_0_1_254), .C2(n_0_152), .ZN(n_0_1_128));
   INV_X1 i_0_1_258 (.A(n_0_1_129), .ZN(n_0_137));
   AOI222_X1 i_0_1_259 (.A1(\temp1[4] [20]), .A2(n_0_1_256), .B1(\temp2[4] [20]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_153), .ZN(n_0_1_129));
   INV_X1 i_0_1_260 (.A(n_0_1_130), .ZN(n_0_138));
   AOI222_X1 i_0_1_261 (.A1(\temp1[4] [21]), .A2(n_0_1_256), .B1(\temp2[4] [21]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_154), .ZN(n_0_1_130));
   INV_X1 i_0_1_262 (.A(n_0_1_131), .ZN(n_0_139));
   AOI222_X1 i_0_1_263 (.A1(\temp1[4] [22]), .A2(n_0_1_256), .B1(\temp2[4] [22]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_155), .ZN(n_0_1_131));
   INV_X1 i_0_1_264 (.A(n_0_1_132), .ZN(n_0_140));
   AOI222_X1 i_0_1_265 (.A1(\temp1[4] [23]), .A2(n_0_1_256), .B1(\temp2[4] [23]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_156), .ZN(n_0_1_132));
   INV_X1 i_0_1_266 (.A(n_0_1_133), .ZN(n_0_141));
   AOI222_X1 i_0_1_267 (.A1(\temp1[4] [24]), .A2(n_0_1_256), .B1(\temp2[4] [24]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_157), .ZN(n_0_1_133));
   INV_X1 i_0_1_268 (.A(n_0_1_134), .ZN(n_0_142));
   AOI222_X1 i_0_1_269 (.A1(\temp1[4] [25]), .A2(n_0_1_256), .B1(\temp2[4] [25]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_158), .ZN(n_0_1_134));
   INV_X1 i_0_1_270 (.A(n_0_1_135), .ZN(n_0_143));
   AOI222_X1 i_0_1_271 (.A1(\temp1[4] [26]), .A2(n_0_1_256), .B1(\temp2[4] [26]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_159), .ZN(n_0_1_135));
   INV_X1 i_0_1_272 (.A(n_0_1_136), .ZN(n_0_144));
   AOI222_X1 i_0_1_273 (.A1(\temp2[4] [27]), .A2(n_0_1_255), .B1(\temp1[4] [27]), 
      .B2(n_0_1_256), .C1(n_0_1_254), .C2(n_0_160), .ZN(n_0_1_136));
   INV_X1 i_0_1_274 (.A(n_0_1_137), .ZN(n_0_145));
   AOI222_X1 i_0_1_275 (.A1(\temp2[4] [28]), .A2(n_0_1_255), .B1(\temp1[4] [28]), 
      .B2(n_0_1_256), .C1(n_0_1_254), .C2(n_0_161), .ZN(n_0_1_137));
   INV_X1 i_0_1_276 (.A(n_0_1_138), .ZN(n_0_146));
   AOI222_X1 i_0_1_277 (.A1(\temp1[4] [29]), .A2(n_0_1_256), .B1(\temp2[4] [29]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_162), .ZN(n_0_1_138));
   INV_X1 i_0_1_278 (.A(n_0_1_139), .ZN(n_0_147));
   AOI222_X1 i_0_1_279 (.A1(\temp1[4] [30]), .A2(n_0_1_256), .B1(\temp2[4] [30]), 
      .B2(n_0_1_255), .C1(n_0_1_254), .C2(n_0_163), .ZN(n_0_1_139));
   INV_X1 i_0_1_280 (.A(n_0_1_140), .ZN(n_0_148));
   AOI221_X1 i_0_1_281 (.A(n_0_1_253), .B1(\temp2[4] [31]), .B2(n_0_1_255), 
      .C1(\temp1[4] [31]), .C2(n_0_1_256), .ZN(n_0_1_140));
   INV_X1 i_0_1_282 (.A(n_0_1_141), .ZN(n_0_150));
   AOI222_X1 i_0_1_283 (.A1(\temp1[3] [18]), .A2(n_0_1_260), .B1(\temp2[3] [18]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_166), .ZN(n_0_1_141));
   INV_X1 i_0_1_284 (.A(n_0_1_142), .ZN(n_0_151));
   AOI222_X1 i_0_1_285 (.A1(\temp1[3] [19]), .A2(n_0_1_260), .B1(\temp2[3] [19]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_167), .ZN(n_0_1_142));
   INV_X1 i_0_1_286 (.A(n_0_1_143), .ZN(n_0_152));
   AOI222_X1 i_0_1_287 (.A1(\temp1[3] [20]), .A2(n_0_1_260), .B1(\temp2[3] [20]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_168), .ZN(n_0_1_143));
   INV_X1 i_0_1_288 (.A(n_0_1_144), .ZN(n_0_153));
   AOI222_X1 i_0_1_289 (.A1(\temp1[3] [21]), .A2(n_0_1_260), .B1(\temp2[3] [21]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_169), .ZN(n_0_1_144));
   INV_X1 i_0_1_290 (.A(n_0_1_145), .ZN(n_0_154));
   AOI222_X1 i_0_1_291 (.A1(\temp1[3] [22]), .A2(n_0_1_260), .B1(\temp2[3] [22]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_170), .ZN(n_0_1_145));
   INV_X1 i_0_1_292 (.A(n_0_1_146), .ZN(n_0_155));
   AOI222_X1 i_0_1_293 (.A1(\temp1[3] [23]), .A2(n_0_1_260), .B1(\temp2[3] [23]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_171), .ZN(n_0_1_146));
   INV_X1 i_0_1_294 (.A(n_0_1_147), .ZN(n_0_156));
   AOI222_X1 i_0_1_295 (.A1(\temp1[3] [24]), .A2(n_0_1_260), .B1(\temp2[3] [24]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_172), .ZN(n_0_1_147));
   INV_X1 i_0_1_296 (.A(n_0_1_148), .ZN(n_0_157));
   AOI222_X1 i_0_1_297 (.A1(\temp1[3] [25]), .A2(n_0_1_260), .B1(\temp2[3] [25]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_173), .ZN(n_0_1_148));
   INV_X1 i_0_1_298 (.A(n_0_1_149), .ZN(n_0_158));
   AOI222_X1 i_0_1_299 (.A1(\temp1[3] [26]), .A2(n_0_1_260), .B1(\temp2[3] [26]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_174), .ZN(n_0_1_149));
   INV_X1 i_0_1_300 (.A(n_0_1_150), .ZN(n_0_159));
   AOI222_X1 i_0_1_301 (.A1(\temp1[3] [27]), .A2(n_0_1_260), .B1(\temp2[3] [27]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_175), .ZN(n_0_1_150));
   INV_X1 i_0_1_302 (.A(n_0_1_151), .ZN(n_0_160));
   AOI222_X1 i_0_1_303 (.A1(\temp1[3] [28]), .A2(n_0_1_260), .B1(\temp2[3] [28]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_176), .ZN(n_0_1_151));
   INV_X1 i_0_1_304 (.A(n_0_1_152), .ZN(n_0_161));
   AOI222_X1 i_0_1_305 (.A1(\temp1[3] [29]), .A2(n_0_1_260), .B1(\temp2[3] [29]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_177), .ZN(n_0_1_152));
   INV_X1 i_0_1_306 (.A(n_0_1_153), .ZN(n_0_162));
   AOI222_X1 i_0_1_307 (.A1(\temp1[3] [30]), .A2(n_0_1_260), .B1(\temp2[3] [30]), 
      .B2(n_0_1_261), .C1(n_0_1_259), .C2(n_0_178), .ZN(n_0_1_153));
   INV_X1 i_0_1_308 (.A(n_0_1_154), .ZN(n_0_163));
   AOI221_X1 i_0_1_309 (.A(n_0_1_258), .B1(\temp2[3] [31]), .B2(n_0_1_261), 
      .C1(\temp1[3] [31]), .C2(n_0_1_260), .ZN(n_0_1_154));
   INV_X1 i_0_1_310 (.A(n_0_1_155), .ZN(n_0_165));
   AOI222_X1 i_0_1_311 (.A1(\temp1[2] [18]), .A2(n_0_1_265), .B1(\temp2[2] [18]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_181), .ZN(n_0_1_155));
   INV_X1 i_0_1_312 (.A(n_0_1_156), .ZN(n_0_166));
   AOI222_X1 i_0_1_313 (.A1(\temp1[2] [19]), .A2(n_0_1_265), .B1(\temp2[2] [19]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_182), .ZN(n_0_1_156));
   INV_X1 i_0_1_314 (.A(n_0_1_157), .ZN(n_0_167));
   AOI222_X1 i_0_1_315 (.A1(\temp1[2] [20]), .A2(n_0_1_265), .B1(\temp2[2] [20]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_183), .ZN(n_0_1_157));
   INV_X1 i_0_1_316 (.A(n_0_1_158), .ZN(n_0_168));
   AOI222_X1 i_0_1_317 (.A1(\temp1[2] [21]), .A2(n_0_1_265), .B1(\temp2[2] [21]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_184), .ZN(n_0_1_158));
   INV_X1 i_0_1_318 (.A(n_0_1_159), .ZN(n_0_169));
   AOI222_X1 i_0_1_319 (.A1(\temp1[2] [22]), .A2(n_0_1_265), .B1(\temp2[2] [22]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_185), .ZN(n_0_1_159));
   INV_X1 i_0_1_320 (.A(n_0_1_160), .ZN(n_0_170));
   AOI222_X1 i_0_1_321 (.A1(\temp1[2] [23]), .A2(n_0_1_265), .B1(\temp2[2] [23]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_186), .ZN(n_0_1_160));
   INV_X1 i_0_1_322 (.A(n_0_1_161), .ZN(n_0_171));
   AOI222_X1 i_0_1_323 (.A1(\temp1[2] [24]), .A2(n_0_1_265), .B1(\temp2[2] [24]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_187), .ZN(n_0_1_161));
   INV_X1 i_0_1_324 (.A(n_0_1_162), .ZN(n_0_172));
   AOI222_X1 i_0_1_325 (.A1(\temp1[2] [25]), .A2(n_0_1_265), .B1(\temp2[2] [25]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_188), .ZN(n_0_1_162));
   INV_X1 i_0_1_326 (.A(n_0_1_163), .ZN(n_0_173));
   AOI222_X1 i_0_1_327 (.A1(\temp1[2] [26]), .A2(n_0_1_265), .B1(\temp2[2] [26]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_189), .ZN(n_0_1_163));
   INV_X1 i_0_1_328 (.A(n_0_1_164), .ZN(n_0_174));
   AOI222_X1 i_0_1_329 (.A1(\temp1[2] [27]), .A2(n_0_1_265), .B1(\temp2[2] [27]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_190), .ZN(n_0_1_164));
   INV_X1 i_0_1_330 (.A(n_0_1_165), .ZN(n_0_175));
   AOI222_X1 i_0_1_331 (.A1(\temp1[2] [28]), .A2(n_0_1_265), .B1(\temp2[2] [28]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_191), .ZN(n_0_1_165));
   INV_X1 i_0_1_332 (.A(n_0_1_166), .ZN(n_0_176));
   AOI222_X1 i_0_1_333 (.A1(\temp1[2] [29]), .A2(n_0_1_265), .B1(\temp2[2] [29]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_192), .ZN(n_0_1_166));
   INV_X1 i_0_1_334 (.A(n_0_1_167), .ZN(n_0_177));
   AOI222_X1 i_0_1_335 (.A1(\temp1[2] [30]), .A2(n_0_1_265), .B1(\temp2[2] [30]), 
      .B2(n_0_1_266), .C1(n_0_1_264), .C2(n_0_193), .ZN(n_0_1_167));
   INV_X1 i_0_1_336 (.A(n_0_1_168), .ZN(n_0_178));
   AOI221_X1 i_0_1_337 (.A(n_0_1_263), .B1(\temp2[2] [31]), .B2(n_0_1_266), 
      .C1(\temp1[2] [31]), .C2(n_0_1_265), .ZN(n_0_1_168));
   INV_X1 i_0_1_338 (.A(n_0_1_169), .ZN(n_0_180));
   AOI222_X1 i_0_1_339 (.A1(r[1]), .A2(n_0_196), .B1(\temp1[1] [18]), .B2(
      n_0_1_268), .C1(\temp2[1] [18]), .C2(n_0_1_271), .ZN(n_0_1_169));
   INV_X1 i_0_1_340 (.A(n_0_1_170), .ZN(n_0_181));
   AOI222_X1 i_0_1_341 (.A1(mn[3]), .A2(n_0_1_270), .B1(\temp1[1] [19]), 
      .B2(n_0_1_268), .C1(\temp2[1] [19]), .C2(n_0_1_271), .ZN(n_0_1_170));
   INV_X1 i_0_1_342 (.A(n_0_1_171), .ZN(n_0_182));
   AOI222_X1 i_0_1_343 (.A1(mn[4]), .A2(n_0_1_270), .B1(\temp1[1] [20]), 
      .B2(n_0_1_268), .C1(\temp2[1] [20]), .C2(n_0_1_271), .ZN(n_0_1_171));
   INV_X1 i_0_1_344 (.A(n_0_1_172), .ZN(n_0_183));
   AOI222_X1 i_0_1_345 (.A1(mn[5]), .A2(n_0_1_270), .B1(\temp1[1] [21]), 
      .B2(n_0_1_268), .C1(\temp2[1] [21]), .C2(n_0_1_271), .ZN(n_0_1_172));
   INV_X1 i_0_1_346 (.A(n_0_1_173), .ZN(n_0_184));
   AOI222_X1 i_0_1_347 (.A1(mn[6]), .A2(n_0_1_270), .B1(\temp1[1] [22]), 
      .B2(n_0_1_268), .C1(\temp2[1] [22]), .C2(n_0_1_271), .ZN(n_0_1_173));
   INV_X1 i_0_1_348 (.A(n_0_1_174), .ZN(n_0_185));
   AOI222_X1 i_0_1_349 (.A1(mn[7]), .A2(n_0_1_270), .B1(\temp1[1] [23]), 
      .B2(n_0_1_268), .C1(\temp2[1] [23]), .C2(n_0_1_271), .ZN(n_0_1_174));
   INV_X1 i_0_1_350 (.A(n_0_1_175), .ZN(n_0_186));
   AOI222_X1 i_0_1_351 (.A1(mn[8]), .A2(n_0_1_270), .B1(\temp1[1] [24]), 
      .B2(n_0_1_268), .C1(\temp2[1] [24]), .C2(n_0_1_271), .ZN(n_0_1_175));
   INV_X1 i_0_1_352 (.A(n_0_1_176), .ZN(n_0_187));
   AOI222_X1 i_0_1_353 (.A1(mn[9]), .A2(n_0_1_270), .B1(\temp1[1] [25]), 
      .B2(n_0_1_268), .C1(\temp2[1] [25]), .C2(n_0_1_271), .ZN(n_0_1_176));
   INV_X1 i_0_1_354 (.A(n_0_1_177), .ZN(n_0_188));
   AOI222_X1 i_0_1_355 (.A1(mn[10]), .A2(n_0_1_270), .B1(\temp1[1] [26]), 
      .B2(n_0_1_268), .C1(\temp2[1] [26]), .C2(n_0_1_271), .ZN(n_0_1_177));
   INV_X1 i_0_1_356 (.A(n_0_1_178), .ZN(n_0_189));
   AOI222_X1 i_0_1_357 (.A1(mn[11]), .A2(n_0_1_270), .B1(\temp1[1] [27]), 
      .B2(n_0_1_268), .C1(\temp2[1] [27]), .C2(n_0_1_271), .ZN(n_0_1_178));
   INV_X1 i_0_1_358 (.A(n_0_1_179), .ZN(n_0_190));
   AOI222_X1 i_0_1_359 (.A1(mn[12]), .A2(n_0_1_270), .B1(\temp1[1] [28]), 
      .B2(n_0_1_268), .C1(\temp2[1] [28]), .C2(n_0_1_271), .ZN(n_0_1_179));
   INV_X1 i_0_1_360 (.A(n_0_1_180), .ZN(n_0_191));
   AOI222_X1 i_0_1_361 (.A1(r[1]), .A2(n_0_207), .B1(\temp1[1] [29]), .B2(
      n_0_1_268), .C1(\temp2[1] [29]), .C2(n_0_1_271), .ZN(n_0_1_180));
   INV_X1 i_0_1_362 (.A(n_0_1_181), .ZN(n_0_192));
   AOI222_X1 i_0_1_363 (.A1(r[1]), .A2(n_0_208), .B1(\temp1[1] [30]), .B2(
      n_0_1_268), .C1(\temp2[1] [30]), .C2(n_0_1_271), .ZN(n_0_1_181));
   INV_X1 i_0_1_364 (.A(n_0_1_182), .ZN(n_0_193));
   AOI221_X1 i_0_1_365 (.A(n_0_1_269), .B1(\temp2[1] [31]), .B2(n_0_1_271), 
      .C1(\temp1[1] [31]), .C2(n_0_1_268), .ZN(n_0_1_182));
   AND2_X1 i_0_1_366 (.A1(r[0]), .A2(mn[1]), .ZN(n_0_195));
   AND2_X1 i_0_1_367 (.A1(r[0]), .A2(mn[2]), .ZN(n_0_196));
   AND2_X1 i_0_1_368 (.A1(r[0]), .A2(mn[3]), .ZN(n_0_197));
   AND2_X1 i_0_1_369 (.A1(r[0]), .A2(mn[4]), .ZN(n_0_198));
   AND2_X1 i_0_1_370 (.A1(r[0]), .A2(mn[5]), .ZN(n_0_199));
   AND2_X1 i_0_1_371 (.A1(r[0]), .A2(mn[6]), .ZN(n_0_200));
   AND2_X1 i_0_1_372 (.A1(r[0]), .A2(mn[7]), .ZN(n_0_201));
   AND2_X1 i_0_1_373 (.A1(r[0]), .A2(mn[8]), .ZN(n_0_202));
   AND2_X1 i_0_1_374 (.A1(r[0]), .A2(mn[9]), .ZN(n_0_203));
   AND2_X1 i_0_1_375 (.A1(r[0]), .A2(mn[10]), .ZN(n_0_204));
   AND2_X1 i_0_1_376 (.A1(r[0]), .A2(mn[11]), .ZN(n_0_205));
   AND2_X1 i_0_1_377 (.A1(r[0]), .A2(mn[12]), .ZN(n_0_206));
   AND2_X1 i_0_1_378 (.A1(r[0]), .A2(mn[13]), .ZN(n_0_207));
   AND2_X1 i_0_1_379 (.A1(r[0]), .A2(mn[14]), .ZN(n_0_208));
   AOI22_X1 i_0_1_380 (.A1(n_0_1_186), .A2(n_0_1_185), .B1(n_0_1_184), .B2(
      n_0_1_183), .ZN(overflow));
   NOR3_X1 i_0_1_381 (.A1(n_0_1_204), .A2(n_0_1_187), .A3(n_0_1_203), .ZN(
      n_0_1_183));
   NOR4_X1 i_0_1_382 (.A1(n_0_1_208), .A2(n_0_1_198), .A3(n_0_1_192), .A4(
      n_0_1_201), .ZN(n_0_1_184));
   AND3_X1 i_0_1_383 (.A1(n_0_1_204), .A2(n_0_1_201), .A3(n_0_1_198), .ZN(
      n_0_1_185));
   AND4_X1 i_0_1_384 (.A1(n_0_1_203), .A2(n_0_1_187), .A3(n_0_1_208), .A4(
      n_0_1_192), .ZN(n_0_1_186));
   AOI222_X1 i_0_1_385 (.A1(\temp2[14] [27]), .A2(n_0_1_276), .B1(
      \temp1[14] [27]), .B2(n_0_1_277), .C1(n_0_1_275), .C2(n_0_10), .ZN(
      n_0_1_187));
   INV_X1 i_0_1_386 (.A(n_0_1_188), .ZN(n_0_10));
   AOI222_X1 i_0_1_387 (.A1(\temp2[13] [28]), .A2(n_0_1_274), .B1(
      \temp1[13] [28]), .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_26), .ZN(
      n_0_1_188));
   INV_X1 i_0_1_388 (.A(n_0_1_189), .ZN(n_0_26));
   AOI222_X1 i_0_1_389 (.A1(\temp2[12] [29]), .A2(n_0_1_215), .B1(
      \temp1[12] [29]), .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_42), .ZN(
      n_0_1_189));
   INV_X1 i_0_1_390 (.A(n_0_1_190), .ZN(n_0_42));
   AOI222_X1 i_0_1_391 (.A1(\temp2[11] [30]), .A2(n_0_1_221), .B1(
      \temp1[11] [30]), .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_58), .ZN(
      n_0_1_190));
   INV_X1 i_0_1_392 (.A(n_0_1_191), .ZN(n_0_58));
   AOI221_X1 i_0_1_393 (.A(n_0_1_223), .B1(\temp2[10] [31]), .B2(n_0_1_226), 
      .C1(\temp1[10] [31]), .C2(n_0_1_225), .ZN(n_0_1_191));
   AOI222_X1 i_0_1_394 (.A1(\temp1[14] [26]), .A2(n_0_1_277), .B1(
      \temp2[14] [26]), .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_9), .ZN(
      n_0_1_192));
   INV_X1 i_0_1_395 (.A(n_0_1_193), .ZN(n_0_9));
   AOI222_X1 i_0_1_396 (.A1(\temp2[13] [27]), .A2(n_0_1_274), .B1(
      \temp1[13] [27]), .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_25), .ZN(
      n_0_1_193));
   INV_X1 i_0_1_397 (.A(n_0_1_194), .ZN(n_0_25));
   AOI222_X1 i_0_1_398 (.A1(\temp2[12] [28]), .A2(n_0_1_215), .B1(
      \temp1[12] [28]), .B2(n_0_1_216), .C1(n_0_1_214), .C2(n_0_41), .ZN(
      n_0_1_194));
   INV_X1 i_0_1_399 (.A(n_0_1_195), .ZN(n_0_41));
   AOI222_X1 i_0_1_400 (.A1(\temp2[11] [29]), .A2(n_0_1_221), .B1(
      \temp1[11] [29]), .B2(n_0_1_220), .C1(n_0_1_219), .C2(n_0_57), .ZN(
      n_0_1_195));
   INV_X1 i_0_1_401 (.A(n_0_1_196), .ZN(n_0_57));
   AOI222_X1 i_0_1_402 (.A1(\temp2[10] [30]), .A2(n_0_1_226), .B1(
      \temp1[10] [30]), .B2(n_0_1_225), .C1(n_0_1_224), .C2(n_0_73), .ZN(
      n_0_1_196));
   INV_X1 i_0_1_403 (.A(n_0_1_197), .ZN(n_0_73));
   AOI221_X1 i_0_1_404 (.A(n_0_1_228), .B1(\temp2[9] [31]), .B2(n_0_1_231), 
      .C1(\temp1[9] [31]), .C2(n_0_1_230), .ZN(n_0_1_197));
   AOI222_X1 i_0_1_405 (.A1(\temp2[14] [29]), .A2(n_0_1_276), .B1(
      \temp1[14] [29]), .B2(n_0_1_277), .C1(n_0_1_275), .C2(n_0_12), .ZN(
      n_0_1_198));
   INV_X1 i_0_1_406 (.A(n_0_1_199), .ZN(n_0_12));
   AOI222_X1 i_0_1_407 (.A1(\temp2[13] [30]), .A2(n_0_1_274), .B1(
      \temp1[13] [30]), .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_28), .ZN(
      n_0_1_199));
   INV_X1 i_0_1_408 (.A(n_0_1_200), .ZN(n_0_28));
   AOI221_X1 i_0_1_409 (.A(n_0_1_213), .B1(\temp2[12] [31]), .B2(n_0_1_215), 
      .C1(\temp1[12] [31]), .C2(n_0_1_216), .ZN(n_0_1_200));
   AOI222_X1 i_0_1_410 (.A1(\temp2[14] [30]), .A2(n_0_1_276), .B1(
      \temp1[14] [30]), .B2(n_0_1_277), .C1(n_0_1_275), .C2(n_0_13), .ZN(
      n_0_1_201));
   INV_X1 i_0_1_411 (.A(n_0_1_202), .ZN(n_0_13));
   AOI221_X1 i_0_1_412 (.A(n_0_1_211), .B1(\temp2[13] [31]), .B2(n_0_1_274), 
      .C1(\temp1[13] [31]), .C2(n_0_1_273), .ZN(n_0_1_202));
   AOI221_X1 i_0_1_413 (.A(n_0_1_209), .B1(\temp2[14] [32]), .B2(n_0_1_276), 
      .C1(\temp1[14] [32]), .C2(n_0_1_277), .ZN(n_0_1_203));
   AOI222_X1 i_0_1_414 (.A1(\temp1[14] [28]), .A2(n_0_1_277), .B1(
      \temp2[14] [28]), .B2(n_0_1_276), .C1(n_0_1_275), .C2(n_0_11), .ZN(
      n_0_1_204));
   INV_X1 i_0_1_415 (.A(n_0_1_205), .ZN(n_0_11));
   AOI222_X1 i_0_1_416 (.A1(\temp2[13] [29]), .A2(n_0_1_274), .B1(
      \temp1[13] [29]), .B2(n_0_1_273), .C1(n_0_1_272), .C2(n_0_27), .ZN(
      n_0_1_205));
   INV_X1 i_0_1_417 (.A(n_0_1_206), .ZN(n_0_27));
   AOI222_X1 i_0_1_418 (.A1(\temp1[12] [30]), .A2(n_0_1_216), .B1(
      \temp2[12] [30]), .B2(n_0_1_215), .C1(n_0_1_214), .C2(n_0_43), .ZN(
      n_0_1_206));
   INV_X1 i_0_1_419 (.A(n_0_1_207), .ZN(n_0_43));
   AOI221_X1 i_0_1_420 (.A(n_0_1_218), .B1(\temp2[11] [31]), .B2(n_0_1_221), 
      .C1(\temp1[11] [31]), .C2(n_0_1_220), .ZN(n_0_1_207));
   AOI221_X1 i_0_1_421 (.A(n_0_1_209), .B1(\temp2[14] [31]), .B2(n_0_1_276), 
      .C1(\temp1[14] [31]), .C2(n_0_1_277), .ZN(n_0_1_208));
   AND2_X1 i_0_1_422 (.A1(n_0_1_275), .A2(n_0_14), .ZN(n_0_1_209));
   INV_X1 i_0_1_423 (.A(n_0_1_210), .ZN(n_0_14));
   AOI221_X1 i_0_1_424 (.A(n_0_1_211), .B1(\temp2[13] [32]), .B2(n_0_1_274), 
      .C1(\temp1[13] [32]), .C2(n_0_1_273), .ZN(n_0_1_210));
   AND2_X1 i_0_1_425 (.A1(n_0_1_272), .A2(n_0_29), .ZN(n_0_1_211));
   INV_X1 i_0_1_426 (.A(n_0_1_212), .ZN(n_0_29));
   AOI221_X1 i_0_1_427 (.A(n_0_1_213), .B1(\temp2[12] [32]), .B2(n_0_1_215), 
      .C1(\temp1[12] [32]), .C2(n_0_1_216), .ZN(n_0_1_212));
   AND2_X1 i_0_1_428 (.A1(n_0_44), .A2(n_0_1_214), .ZN(n_0_1_213));
   NOR2_X1 i_0_1_429 (.A1(n_0_1_216), .A2(n_0_1_215), .ZN(n_0_1_214));
   NOR2_X1 i_0_1_430 (.A1(n_0_1_289), .A2(r[11]), .ZN(n_0_1_215));
   NOR2_X1 i_0_1_431 (.A1(r[12]), .A2(n_0_1_288), .ZN(n_0_1_216));
   INV_X1 i_0_1_432 (.A(n_0_1_217), .ZN(n_0_44));
   AOI221_X1 i_0_1_433 (.A(n_0_1_218), .B1(\temp2[11] [32]), .B2(n_0_1_221), 
      .C1(\temp1[11] [32]), .C2(n_0_1_220), .ZN(n_0_1_217));
   AND2_X1 i_0_1_434 (.A1(n_0_59), .A2(n_0_1_219), .ZN(n_0_1_218));
   NOR2_X1 i_0_1_435 (.A1(n_0_1_221), .A2(n_0_1_220), .ZN(n_0_1_219));
   NOR2_X1 i_0_1_436 (.A1(r[11]), .A2(n_0_1_287), .ZN(n_0_1_220));
   NOR2_X1 i_0_1_437 (.A1(n_0_1_288), .A2(r[10]), .ZN(n_0_1_221));
   INV_X1 i_0_1_438 (.A(n_0_1_222), .ZN(n_0_59));
   AOI221_X1 i_0_1_439 (.A(n_0_1_223), .B1(\temp2[10] [32]), .B2(n_0_1_226), 
      .C1(\temp1[10] [32]), .C2(n_0_1_225), .ZN(n_0_1_222));
   AND2_X1 i_0_1_440 (.A1(n_0_74), .A2(n_0_1_224), .ZN(n_0_1_223));
   NOR2_X1 i_0_1_441 (.A1(n_0_1_226), .A2(n_0_1_225), .ZN(n_0_1_224));
   NOR2_X1 i_0_1_442 (.A1(r[10]), .A2(n_0_1_286), .ZN(n_0_1_225));
   NOR2_X1 i_0_1_443 (.A1(n_0_1_287), .A2(r[9]), .ZN(n_0_1_226));
   INV_X1 i_0_1_444 (.A(n_0_1_227), .ZN(n_0_74));
   AOI221_X1 i_0_1_445 (.A(n_0_1_228), .B1(\temp2[9] [32]), .B2(n_0_1_231), 
      .C1(\temp1[9] [32]), .C2(n_0_1_230), .ZN(n_0_1_227));
   AND2_X1 i_0_1_446 (.A1(n_0_89), .A2(n_0_1_229), .ZN(n_0_1_228));
   NOR2_X1 i_0_1_447 (.A1(n_0_1_231), .A2(n_0_1_230), .ZN(n_0_1_229));
   NOR2_X1 i_0_1_448 (.A1(r[9]), .A2(n_0_1_285), .ZN(n_0_1_230));
   NOR2_X1 i_0_1_449 (.A1(n_0_1_286), .A2(r[8]), .ZN(n_0_1_231));
   INV_X1 i_0_1_450 (.A(n_0_1_232), .ZN(n_0_89));
   AOI221_X1 i_0_1_451 (.A(n_0_1_233), .B1(\temp2[8] [32]), .B2(n_0_1_236), 
      .C1(\temp1[8] [32]), .C2(n_0_1_235), .ZN(n_0_1_232));
   AND2_X1 i_0_1_452 (.A1(n_0_104), .A2(n_0_1_234), .ZN(n_0_1_233));
   NOR2_X1 i_0_1_453 (.A1(n_0_1_236), .A2(n_0_1_235), .ZN(n_0_1_234));
   NOR2_X1 i_0_1_454 (.A1(r[8]), .A2(n_0_1_284), .ZN(n_0_1_235));
   NOR2_X1 i_0_1_455 (.A1(n_0_1_285), .A2(r[7]), .ZN(n_0_1_236));
   INV_X1 i_0_1_456 (.A(n_0_1_237), .ZN(n_0_104));
   AOI221_X1 i_0_1_457 (.A(n_0_1_238), .B1(\temp2[7] [32]), .B2(n_0_1_240), 
      .C1(\temp1[7] [32]), .C2(n_0_1_241), .ZN(n_0_1_237));
   AND2_X1 i_0_1_458 (.A1(n_0_119), .A2(n_0_1_239), .ZN(n_0_1_238));
   NOR2_X1 i_0_1_459 (.A1(n_0_1_241), .A2(n_0_1_240), .ZN(n_0_1_239));
   NOR2_X1 i_0_1_460 (.A1(n_0_1_284), .A2(r[6]), .ZN(n_0_1_240));
   NOR2_X1 i_0_1_461 (.A1(r[7]), .A2(n_0_1_283), .ZN(n_0_1_241));
   INV_X1 i_0_1_462 (.A(n_0_1_242), .ZN(n_0_119));
   AOI221_X1 i_0_1_463 (.A(n_0_1_243), .B1(\temp2[6] [32]), .B2(n_0_1_246), 
      .C1(\temp1[6] [32]), .C2(n_0_1_245), .ZN(n_0_1_242));
   AND2_X1 i_0_1_464 (.A1(n_0_134), .A2(n_0_1_244), .ZN(n_0_1_243));
   NOR2_X1 i_0_1_465 (.A1(n_0_1_246), .A2(n_0_1_245), .ZN(n_0_1_244));
   NOR2_X1 i_0_1_466 (.A1(r[6]), .A2(n_0_1_282), .ZN(n_0_1_245));
   NOR2_X1 i_0_1_467 (.A1(n_0_1_283), .A2(r[5]), .ZN(n_0_1_246));
   INV_X1 i_0_1_468 (.A(n_0_1_247), .ZN(n_0_134));
   AOI221_X1 i_0_1_469 (.A(n_0_1_248), .B1(\temp2[5] [32]), .B2(n_0_1_251), 
      .C1(\temp1[5] [32]), .C2(n_0_1_250), .ZN(n_0_1_247));
   AND2_X1 i_0_1_470 (.A1(n_0_149), .A2(n_0_1_249), .ZN(n_0_1_248));
   NOR2_X1 i_0_1_471 (.A1(n_0_1_251), .A2(n_0_1_250), .ZN(n_0_1_249));
   NOR2_X1 i_0_1_472 (.A1(r[5]), .A2(n_0_1_281), .ZN(n_0_1_250));
   NOR2_X1 i_0_1_473 (.A1(n_0_1_282), .A2(r[4]), .ZN(n_0_1_251));
   INV_X1 i_0_1_474 (.A(n_0_1_252), .ZN(n_0_149));
   AOI221_X1 i_0_1_475 (.A(n_0_1_253), .B1(\temp2[4] [32]), .B2(n_0_1_255), 
      .C1(\temp1[4] [32]), .C2(n_0_1_256), .ZN(n_0_1_252));
   AND2_X1 i_0_1_476 (.A1(n_0_164), .A2(n_0_1_254), .ZN(n_0_1_253));
   NOR2_X1 i_0_1_477 (.A1(n_0_1_256), .A2(n_0_1_255), .ZN(n_0_1_254));
   NOR2_X1 i_0_1_478 (.A1(n_0_1_281), .A2(r[3]), .ZN(n_0_1_255));
   NOR2_X1 i_0_1_479 (.A1(r[4]), .A2(n_0_1_280), .ZN(n_0_1_256));
   INV_X1 i_0_1_480 (.A(n_0_1_257), .ZN(n_0_164));
   AOI221_X1 i_0_1_481 (.A(n_0_1_258), .B1(\temp2[3] [32]), .B2(n_0_1_261), 
      .C1(\temp1[3] [32]), .C2(n_0_1_260), .ZN(n_0_1_257));
   AND2_X1 i_0_1_482 (.A1(n_0_179), .A2(n_0_1_259), .ZN(n_0_1_258));
   NOR2_X1 i_0_1_483 (.A1(n_0_1_261), .A2(n_0_1_260), .ZN(n_0_1_259));
   NOR2_X1 i_0_1_484 (.A1(r[3]), .A2(n_0_1_279), .ZN(n_0_1_260));
   NOR2_X1 i_0_1_485 (.A1(n_0_1_280), .A2(r[2]), .ZN(n_0_1_261));
   INV_X1 i_0_1_486 (.A(n_0_1_262), .ZN(n_0_179));
   AOI221_X1 i_0_1_487 (.A(n_0_1_263), .B1(\temp2[2] [32]), .B2(n_0_1_266), 
      .C1(\temp1[2] [32]), .C2(n_0_1_265), .ZN(n_0_1_262));
   AND2_X1 i_0_1_488 (.A1(n_0_194), .A2(n_0_1_264), .ZN(n_0_1_263));
   NOR2_X1 i_0_1_489 (.A1(n_0_1_266), .A2(n_0_1_265), .ZN(n_0_1_264));
   NOR2_X1 i_0_1_490 (.A1(r[2]), .A2(n_0_1_278), .ZN(n_0_1_265));
   NOR2_X1 i_0_1_491 (.A1(n_0_1_279), .A2(r[1]), .ZN(n_0_1_266));
   INV_X1 i_0_1_492 (.A(n_0_1_267), .ZN(n_0_194));
   AOI221_X1 i_0_1_493 (.A(n_0_1_269), .B1(\temp1[1] [32]), .B2(n_0_1_268), 
      .C1(\temp2[1] [32]), .C2(n_0_1_271), .ZN(n_0_1_267));
   AND2_X1 i_0_1_494 (.A1(n_0_1_278), .A2(r[0]), .ZN(n_0_1_268));
   AND2_X1 i_0_1_495 (.A1(r[1]), .A2(n_0_209), .ZN(n_0_1_269));
   AND2_X1 i_0_1_496 (.A1(r[1]), .A2(r[0]), .ZN(n_0_1_270));
   AND2_X1 i_0_1_497 (.A1(r[0]), .A2(mn[15]), .ZN(n_0_209));
   NOR2_X1 i_0_1_498 (.A1(n_0_1_278), .A2(r[0]), .ZN(n_0_1_271));
   NOR2_X1 i_0_1_499 (.A1(n_0_1_274), .A2(n_0_1_273), .ZN(n_0_1_272));
   NOR2_X1 i_0_1_500 (.A1(r[13]), .A2(n_0_1_289), .ZN(n_0_1_273));
   NOR2_X1 i_0_1_501 (.A1(n_0_1_290), .A2(r[12]), .ZN(n_0_1_274));
   NOR2_X1 i_0_1_502 (.A1(n_0_1_277), .A2(n_0_1_276), .ZN(n_0_1_275));
   AND2_X1 i_0_1_503 (.A1(r[14]), .A2(n_0_1_290), .ZN(n_0_1_276));
   NOR2_X1 i_0_1_504 (.A1(r[14]), .A2(n_0_1_290), .ZN(n_0_1_277));
   INV_X1 i_0_1_505 (.A(r[1]), .ZN(n_0_1_278));
   INV_X1 i_0_1_506 (.A(r[2]), .ZN(n_0_1_279));
   INV_X1 i_0_1_507 (.A(r[3]), .ZN(n_0_1_280));
   INV_X1 i_0_1_508 (.A(r[4]), .ZN(n_0_1_281));
   INV_X1 i_0_1_509 (.A(r[5]), .ZN(n_0_1_282));
   INV_X1 i_0_1_510 (.A(r[6]), .ZN(n_0_1_283));
   INV_X1 i_0_1_511 (.A(r[7]), .ZN(n_0_1_284));
   INV_X1 i_0_1_512 (.A(r[8]), .ZN(n_0_1_285));
   INV_X1 i_0_1_513 (.A(r[9]), .ZN(n_0_1_286));
   INV_X1 i_0_1_514 (.A(r[10]), .ZN(n_0_1_287));
   INV_X1 i_0_1_515 (.A(r[11]), .ZN(n_0_1_288));
   INV_X1 i_0_1_516 (.A(r[12]), .ZN(n_0_1_289));
   INV_X1 i_0_1_517 (.A(r[13]), .ZN(n_0_1_290));
endmodule
