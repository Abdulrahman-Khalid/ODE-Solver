/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 18:24:34 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2181230635 */

module Partial_Full_Adder__0_234(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(B), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_230(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_226(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_222(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_218(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_214(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_210(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_206(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_202(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_198(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_194(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_190(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_186(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_182(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_178(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_174(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(S));
   AND2_X1 i_0_1 (.A1(A), .A2(B), .ZN(G));
endmodule

module Carry_Look_Ahead_generic__0_326(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;

   Partial_Full_Adder__0_234 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(), .B(B[16]), 
      .Cin(n_29), .S(S[16]), .P(), .G());
   Partial_Full_Adder__0_230 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_30), .S(S[15]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_226 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_31), .S(S[14]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_222 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_32), .S(S[13]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_218 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_33), .S(S[12]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_214 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_34), .S(S[11]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_210 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_35), .S(S[10]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_206 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_36), .S(S[9]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_202 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_37), .S(S[8]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_198 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), 
      .B(B[7]), .Cin(n_38), .S(S[7]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_194 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), 
      .B(B[6]), .Cin(n_39), .S(S[6]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_190 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), 
      .B(B[5]), .Cin(n_40), .S(S[5]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_186 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), 
      .B(B[4]), .Cin(n_41), .S(S[4]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_182 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), 
      .B(B[3]), .Cin(n_42), .S(S[3]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_178 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), 
      .B(B[2]), .Cin(n_28), .S(S[2]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_174 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), 
      .B(B[1]), .Cin(), .S(S[1]), .P(), .G(n_28));
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   AND2_X1 i_1_0 (.A1(B[16]), .A2(n_29), .ZN(S[17]));
   INV_X1 i_1_1 (.A(n_1_0), .ZN(n_29));
   AOI21_X1 i_1_2 (.A(n_0), .B1(n_1), .B2(n_30), .ZN(n_1_0));
   INV_X1 i_1_3 (.A(n_1_1), .ZN(n_30));
   AOI21_X1 i_1_4 (.A(n_2), .B1(n_3), .B2(n_31), .ZN(n_1_1));
   INV_X1 i_1_5 (.A(n_1_2), .ZN(n_31));
   AOI21_X1 i_1_6 (.A(n_4), .B1(n_5), .B2(n_32), .ZN(n_1_2));
   INV_X1 i_1_7 (.A(n_1_3), .ZN(n_32));
   AOI21_X1 i_1_8 (.A(n_6), .B1(n_7), .B2(n_33), .ZN(n_1_3));
   INV_X1 i_1_9 (.A(n_1_4), .ZN(n_33));
   AOI21_X1 i_1_10 (.A(n_8), .B1(n_9), .B2(n_34), .ZN(n_1_4));
   INV_X1 i_1_11 (.A(n_1_5), .ZN(n_34));
   AOI21_X1 i_1_12 (.A(n_10), .B1(n_11), .B2(n_35), .ZN(n_1_5));
   INV_X1 i_1_13 (.A(n_1_6), .ZN(n_35));
   AOI21_X1 i_1_14 (.A(n_12), .B1(n_13), .B2(n_36), .ZN(n_1_6));
   INV_X1 i_1_15 (.A(n_1_7), .ZN(n_36));
   AOI21_X1 i_1_16 (.A(n_14), .B1(n_15), .B2(n_37), .ZN(n_1_7));
   INV_X1 i_1_17 (.A(n_1_8), .ZN(n_37));
   AOI21_X1 i_1_18 (.A(n_16), .B1(n_17), .B2(n_38), .ZN(n_1_8));
   INV_X1 i_1_19 (.A(n_1_9), .ZN(n_38));
   AOI21_X1 i_1_20 (.A(n_18), .B1(n_19), .B2(n_39), .ZN(n_1_9));
   INV_X1 i_1_21 (.A(n_1_10), .ZN(n_39));
   AOI21_X1 i_1_22 (.A(n_20), .B1(n_21), .B2(n_40), .ZN(n_1_10));
   INV_X1 i_1_23 (.A(n_1_11), .ZN(n_40));
   AOI21_X1 i_1_24 (.A(n_22), .B1(n_23), .B2(n_41), .ZN(n_1_11));
   INV_X1 i_1_25 (.A(n_1_12), .ZN(n_41));
   AOI21_X1 i_1_26 (.A(n_24), .B1(n_25), .B2(n_42), .ZN(n_1_12));
   INV_X1 i_1_27 (.A(n_1_13), .ZN(n_42));
   AOI21_X1 i_1_28 (.A(n_26), .B1(n_28), .B2(n_27), .ZN(n_1_13));
endmodule

module MuxCustom__0_2447(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
   AND2_X1 i_0_24 (.A1(selector), .A2(A[24]), .ZN(Y[24]));
   AND2_X1 i_0_25 (.A1(selector), .A2(A[25]), .ZN(Y[25]));
   AND2_X1 i_0_26 (.A1(selector), .A2(A[26]), .ZN(Y[26]));
   AND2_X1 i_0_27 (.A1(selector), .A2(A[27]), .ZN(Y[27]));
   AND2_X1 i_0_28 (.A1(selector), .A2(A[28]), .ZN(Y[28]));
   AND2_X1 i_0_29 (.A1(selector), .A2(A[29]), .ZN(Y[29]));
   AND2_X1 i_0_30 (.A1(selector), .A2(A[30]), .ZN(Y[30]));
endmodule

module MuxCustom__0_2449(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
   AND2_X1 i_0_24 (.A1(selector), .A2(A[24]), .ZN(Y[24]));
   AND2_X1 i_0_25 (.A1(selector), .A2(A[25]), .ZN(Y[25]));
   AND2_X1 i_0_26 (.A1(selector), .A2(A[26]), .ZN(Y[26]));
   AND2_X1 i_0_27 (.A1(selector), .A2(A[27]), .ZN(Y[27]));
   AND2_X1 i_0_28 (.A1(selector), .A2(A[28]), .ZN(Y[28]));
   AND2_X1 i_0_29 (.A1(selector), .A2(A[29]), .ZN(Y[29]));
endmodule

module MuxCustom__0_2451(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
   AND2_X1 i_0_24 (.A1(selector), .A2(A[24]), .ZN(Y[24]));
   AND2_X1 i_0_25 (.A1(selector), .A2(A[25]), .ZN(Y[25]));
   AND2_X1 i_0_26 (.A1(selector), .A2(A[26]), .ZN(Y[26]));
   AND2_X1 i_0_27 (.A1(selector), .A2(A[27]), .ZN(Y[27]));
   AND2_X1 i_0_28 (.A1(selector), .A2(A[28]), .ZN(Y[28]));
endmodule

module MuxCustom__0_2453(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
   AND2_X1 i_0_24 (.A1(selector), .A2(A[24]), .ZN(Y[24]));
   AND2_X1 i_0_25 (.A1(selector), .A2(A[25]), .ZN(Y[25]));
   AND2_X1 i_0_26 (.A1(selector), .A2(A[26]), .ZN(Y[26]));
   AND2_X1 i_0_27 (.A1(selector), .A2(A[27]), .ZN(Y[27]));
endmodule

module MuxCustom__0_2455(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
   AND2_X1 i_0_24 (.A1(selector), .A2(A[24]), .ZN(Y[24]));
   AND2_X1 i_0_25 (.A1(selector), .A2(A[25]), .ZN(Y[25]));
   AND2_X1 i_0_26 (.A1(selector), .A2(A[26]), .ZN(Y[26]));
endmodule

module MuxCustom__0_2457(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
   AND2_X1 i_0_24 (.A1(selector), .A2(A[24]), .ZN(Y[24]));
   AND2_X1 i_0_25 (.A1(selector), .A2(A[25]), .ZN(Y[25]));
endmodule

module MuxCustom__0_2459(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
   AND2_X1 i_0_24 (.A1(selector), .A2(A[24]), .ZN(Y[24]));
endmodule

module MuxCustom__0_2461(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
   AND2_X1 i_0_23 (.A1(selector), .A2(A[23]), .ZN(Y[23]));
endmodule

module MuxCustom__0_2463(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
   AND2_X1 i_0_22 (.A1(selector), .A2(A[22]), .ZN(Y[22]));
endmodule

module MuxCustom__0_2465(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_6 (.A1(selector), .A2(A[6]), .ZN(Y[6]));
   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
   AND2_X1 i_0_21 (.A1(selector), .A2(A[21]), .ZN(Y[21]));
endmodule

module MuxCustom__0_2467(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_5 (.A1(selector), .A2(A[5]), .ZN(Y[5]));
   AND2_X1 i_0_6 (.A1(selector), .A2(A[6]), .ZN(Y[6]));
   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
   AND2_X1 i_0_20 (.A1(selector), .A2(A[20]), .ZN(Y[20]));
endmodule

module MuxCustom__0_2469(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_4 (.A1(selector), .A2(A[4]), .ZN(Y[4]));
   AND2_X1 i_0_5 (.A1(selector), .A2(A[5]), .ZN(Y[5]));
   AND2_X1 i_0_6 (.A1(selector), .A2(A[6]), .ZN(Y[6]));
   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
   AND2_X1 i_0_19 (.A1(selector), .A2(A[19]), .ZN(Y[19]));
endmodule

module MuxCustom__0_2471(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_3 (.A1(selector), .A2(A[3]), .ZN(Y[3]));
   AND2_X1 i_0_4 (.A1(selector), .A2(A[4]), .ZN(Y[4]));
   AND2_X1 i_0_5 (.A1(selector), .A2(A[5]), .ZN(Y[5]));
   AND2_X1 i_0_6 (.A1(selector), .A2(A[6]), .ZN(Y[6]));
   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
   AND2_X1 i_0_18 (.A1(selector), .A2(A[18]), .ZN(Y[18]));
endmodule

module MuxCustom__0_2473(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_2 (.A1(selector), .A2(A[2]), .ZN(Y[2]));
   AND2_X1 i_0_3 (.A1(selector), .A2(A[3]), .ZN(Y[3]));
   AND2_X1 i_0_4 (.A1(selector), .A2(A[4]), .ZN(Y[4]));
   AND2_X1 i_0_5 (.A1(selector), .A2(A[5]), .ZN(Y[5]));
   AND2_X1 i_0_6 (.A1(selector), .A2(A[6]), .ZN(Y[6]));
   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
   AND2_X1 i_0_17 (.A1(selector), .A2(A[17]), .ZN(Y[17]));
endmodule

module MuxCustom__0_2475(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_1 (.A1(selector), .A2(A[1]), .ZN(Y[1]));
   AND2_X1 i_0_2 (.A1(selector), .A2(A[2]), .ZN(Y[2]));
   AND2_X1 i_0_3 (.A1(selector), .A2(A[3]), .ZN(Y[3]));
   AND2_X1 i_0_4 (.A1(selector), .A2(A[4]), .ZN(Y[4]));
   AND2_X1 i_0_5 (.A1(selector), .A2(A[5]), .ZN(Y[5]));
   AND2_X1 i_0_6 (.A1(selector), .A2(A[6]), .ZN(Y[6]));
   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
   AND2_X1 i_0_16 (.A1(selector), .A2(A[16]), .ZN(Y[16]));
endmodule

module MuxCustom(A, Y, selector);
   input [31:0]A;
   output [31:0]Y;
   input selector;

   AND2_X1 i_0_0 (.A1(A[0]), .A2(selector), .ZN(Y[0]));
   AND2_X1 i_0_1 (.A1(selector), .A2(A[1]), .ZN(Y[1]));
   AND2_X1 i_0_2 (.A1(selector), .A2(A[2]), .ZN(Y[2]));
   AND2_X1 i_0_3 (.A1(selector), .A2(A[3]), .ZN(Y[3]));
   AND2_X1 i_0_4 (.A1(selector), .A2(A[4]), .ZN(Y[4]));
   AND2_X1 i_0_5 (.A1(selector), .A2(A[5]), .ZN(Y[5]));
   AND2_X1 i_0_6 (.A1(selector), .A2(A[6]), .ZN(Y[6]));
   AND2_X1 i_0_7 (.A1(selector), .A2(A[7]), .ZN(Y[7]));
   AND2_X1 i_0_8 (.A1(selector), .A2(A[8]), .ZN(Y[8]));
   AND2_X1 i_0_9 (.A1(selector), .A2(A[9]), .ZN(Y[9]));
   AND2_X1 i_0_10 (.A1(selector), .A2(A[10]), .ZN(Y[10]));
   AND2_X1 i_0_11 (.A1(selector), .A2(A[11]), .ZN(Y[11]));
   AND2_X1 i_0_12 (.A1(selector), .A2(A[12]), .ZN(Y[12]));
   AND2_X1 i_0_13 (.A1(selector), .A2(A[13]), .ZN(Y[13]));
   AND2_X1 i_0_14 (.A1(selector), .A2(A[14]), .ZN(Y[14]));
   AND2_X1 i_0_15 (.A1(selector), .A2(A[15]), .ZN(Y[15]));
endmodule

module Partial_Full_Adder__0_401(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_397(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_393(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_389(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_385(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_381(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_377(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_373(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_369(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_365(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_361(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_357(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_353(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_349(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_345(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_341(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_337(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_333(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_489(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_401 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_32), .S(S[17]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_397 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_33), .S(S[16]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_393 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_34), .S(S[15]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_389 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_35), .S(S[14]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_385 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_36), .S(S[13]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_381 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_37), .S(S[12]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_377 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_38), .S(S[11]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_373 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_39), .S(S[10]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_369 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_40), .S(S[9]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_365 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_41), .S(S[8]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_361 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), 
      .B(B[7]), .Cin(n_42), .S(S[7]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_357 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), 
      .B(B[6]), .Cin(n_43), .S(S[6]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_353 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), 
      .B(B[5]), .Cin(n_44), .S(S[5]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_349 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), 
      .B(B[4]), .Cin(n_45), .S(S[4]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_345 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), 
      .B(B[3]), .Cin(n_46), .S(S[3]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_341 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), 
      .B(B[2]), .Cin(n_47), .S(S[2]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_337 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_48), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_333 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[18]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[1]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(Cin), .A2(A[0]), .ZN(n_48));
endmodule

module Partial_Full_Adder__0_568(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_564(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_560(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_556(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_552(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_548(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_544(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_540(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_536(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_532(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_528(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_524(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_520(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_516(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_512(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_508(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_504(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_500(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_496(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_652(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_568 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_32), .S(S[18]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_564 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_33), .S(S[17]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_560 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_34), .S(S[16]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_556 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_35), .S(S[15]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_552 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_36), .S(S[14]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_548 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_37), .S(S[13]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_544 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_38), .S(S[12]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_540 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_39), .S(S[11]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_536 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_40), .S(S[10]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_532 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_41), .S(S[9]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_528 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_42), .S(S[8]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_524 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), 
      .B(B[7]), .Cin(n_43), .S(S[7]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_520 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), 
      .B(B[6]), .Cin(n_44), .S(S[6]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_516 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), 
      .B(B[5]), .Cin(n_45), .S(S[5]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_512 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), 
      .B(B[4]), .Cin(n_46), .S(S[4]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_508 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), 
      .B(B[3]), .Cin(n_47), .S(S[3]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_504 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_48), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_500 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_49), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_496 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[19]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[2]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[1]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(Cin), .A2(A[0]), .ZN(n_49));
endmodule

module Partial_Full_Adder__0_735(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_731(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_727(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_723(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_719(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_715(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_711(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_707(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_703(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_699(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_695(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_691(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_687(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_683(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_679(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_675(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_671(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_667(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_663(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_659(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_815(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_735 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_32), .S(S[19]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_731 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_33), .S(S[18]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_727 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_34), .S(S[17]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_723 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_35), .S(S[16]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_719 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_36), .S(S[15]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_715 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_37), .S(S[14]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_711 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_38), .S(S[13]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_707 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_39), .S(S[12]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_703 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_40), .S(S[11]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_699 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_41), .S(S[10]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_695 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_42), .S(S[9]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_691 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_43), .S(S[8]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_687 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), 
      .B(B[7]), .Cin(n_44), .S(S[7]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_683 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), 
      .B(B[6]), .Cin(n_45), .S(S[6]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_679 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), 
      .B(B[5]), .Cin(n_46), .S(S[5]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_675 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), 
      .B(B[4]), .Cin(n_47), .S(S[4]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_671 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_48), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_667 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_49), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_663 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_50), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_659 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[20]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[3]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[2]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[1]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(Cin), .A2(A[0]), .ZN(n_50));
endmodule

module Partial_Full_Adder__0_902(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_898(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_894(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_890(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_886(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_882(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_878(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_874(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_870(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_866(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_862(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_858(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_854(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_850(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_846(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_842(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_838(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_834(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_830(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_826(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_822(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_978(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_902 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_32), .S(S[20]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_898 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_33), .S(S[19]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_894 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_34), .S(S[18]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_890 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_35), .S(S[17]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_886 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_36), .S(S[16]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_882 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_37), .S(S[15]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_878 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_38), .S(S[14]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_874 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_39), .S(S[13]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_870 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_40), .S(S[12]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_866 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_41), .S(S[11]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_862 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_42), .S(S[10]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_858 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_43), .S(S[9]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_854 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_44), .S(S[8]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_850 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), 
      .B(B[7]), .Cin(n_45), .S(S[7]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_846 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), 
      .B(B[6]), .Cin(n_46), .S(S[6]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_842 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), 
      .B(B[5]), .Cin(n_47), .S(S[5]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_838 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_48), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_834 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_49), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_830 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_50), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_826 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_51), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_822 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[21]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[4]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[3]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[2]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[1]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(Cin), .A2(A[0]), .ZN(n_51));
endmodule

module Partial_Full_Adder__0_1069(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1065(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1061(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1057(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1053(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1049(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1045(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1041(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1037(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1033(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1029(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1025(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1021(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1017(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1013(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1009(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1005(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1001(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_997(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_993(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_989(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_985(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_1141(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_1069 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_32), .S(S[21]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1065 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_33), .S(S[20]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1061 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_34), .S(S[19]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1057 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_35), .S(S[18]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1053 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_36), .S(S[17]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1049 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_37), .S(S[16]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1045 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_38), .S(S[15]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1041 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_39), .S(S[14]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1037 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_40), .S(S[13]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1033 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_41), .S(S[12]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1029 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_42), .S(S[11]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1025 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_43), .S(S[10]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1021 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_44), .S(S[9]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1017 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_45), .S(S[8]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_1013 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), 
      .B(B[7]), .Cin(n_46), .S(S[7]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_1009 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), 
      .B(B[6]), .Cin(n_47), .S(S[6]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_1005 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_48), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_1001 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_49), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_997 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_50), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_993 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_51), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_989 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_52), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_985 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[22]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[5]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[4]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[3]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[2]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[1]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(Cin), .A2(A[0]), .ZN(n_52));
endmodule

module Partial_Full_Adder__0_1236(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1232(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1228(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1224(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1220(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1216(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1212(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1208(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1204(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1200(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1196(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1192(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1188(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1184(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1180(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1176(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1172(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1168(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1164(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1160(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1156(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1152(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1148(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_1304(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_1236 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_32), .S(S[22]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1232 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_33), .S(S[21]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1228 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_34), .S(S[20]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1224 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_35), .S(S[19]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1220 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_36), .S(S[18]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1216 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_37), .S(S[17]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1212 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_38), .S(S[16]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1208 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_39), .S(S[15]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1204 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_40), .S(S[14]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1200 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_41), .S(S[13]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1196 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_42), .S(S[12]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1192 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_43), .S(S[11]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1188 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_44), .S(S[10]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1184 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_45), .S(S[9]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_1180 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_46), .S(S[8]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_1176 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), 
      .B(B[7]), .Cin(n_47), .S(S[7]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_1172 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_48), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_1168 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_49), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_1164 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_50), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_1160 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_51), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_1156 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_52), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_1152 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_53), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_1148 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[23]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[6]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[5]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[4]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[3]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[2]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[1]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(Cin), .A2(A[0]), .ZN(n_53));
endmodule

module Partial_Full_Adder__0_1403(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1399(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1395(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1391(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1387(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1383(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1379(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1375(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1371(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1367(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1363(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1359(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1355(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1351(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1347(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1343(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1339(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1335(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1331(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1327(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1323(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1319(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1315(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1311(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_1467(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_1403 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_32), .S(S[23]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1399 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_33), .S(S[22]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1395 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_34), .S(S[21]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1391 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_35), .S(S[20]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1387 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_36), .S(S[19]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1383 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_37), .S(S[18]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1379 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_38), .S(S[17]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1375 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_39), .S(S[16]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1371 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_40), .S(S[15]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1367 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_41), .S(S[14]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1363 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_42), .S(S[13]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1359 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_43), .S(S[12]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1355 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_44), .S(S[11]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1351 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_45), .S(S[10]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_1347 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_46), .S(S[9]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_1343 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), 
      .B(B[8]), .Cin(n_47), .S(S[8]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_1339 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_48), .S(S[7]), .P(), .G());
   Partial_Full_Adder__0_1335 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_49), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_1331 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_50), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_1327 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_51), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_1323 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_52), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_1319 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_53), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_1315 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_54), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_1311 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[24]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[7]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[6]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[5]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[4]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[3]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[2]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(A[1]), .A2(n_54), .ZN(n_53));
   AND2_X1 i_1_39 (.A1(Cin), .A2(A[0]), .ZN(n_54));
endmodule

module Partial_Full_Adder__0_1570(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1566(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1562(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1558(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1554(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1550(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1546(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1542(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1538(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1534(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1530(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1526(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1522(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1518(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1514(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1510(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1506(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1502(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1498(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1494(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1490(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1486(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1482(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1478(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1474(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_1630(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_1570 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_32), .S(S[24]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1566 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_33), .S(S[23]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1562 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_34), .S(S[22]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1558 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_35), .S(S[21]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1554 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_36), .S(S[20]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1550 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_37), .S(S[19]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1546 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_38), .S(S[18]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1542 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_39), .S(S[17]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1538 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_40), .S(S[16]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1534 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_41), .S(S[15]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1530 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_42), .S(S[14]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1526 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_43), .S(S[13]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1522 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_44), .S(S[12]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1518 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_45), .S(S[11]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_1514 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_46), .S(S[10]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_1510 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), 
      .B(B[9]), .Cin(n_47), .S(S[9]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_1506 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), .B(), 
      .Cin(n_48), .S(S[8]), .P(), .G());
   Partial_Full_Adder__0_1502 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_49), .S(S[7]), .P(), .G());
   Partial_Full_Adder__0_1498 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_50), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_1494 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_51), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_1490 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_52), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_1486 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_53), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_1482 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_54), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_1478 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_55), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_1474 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[25]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[8]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[7]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[6]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[5]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[4]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[3]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(A[2]), .A2(n_54), .ZN(n_53));
   AND2_X1 i_1_39 (.A1(A[1]), .A2(n_55), .ZN(n_54));
   AND2_X1 i_1_40 (.A1(Cin), .A2(A[0]), .ZN(n_55));
endmodule

module Partial_Full_Adder__0_1737(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1733(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1729(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1725(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1721(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1717(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1713(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1709(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1705(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1701(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1697(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1693(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1689(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1685(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1681(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1677(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1673(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1669(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1665(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1661(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1657(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1653(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1649(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1645(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1641(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1637(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_1793(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_1737 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_32), .S(S[25]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1733 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_33), .S(S[24]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1729 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_34), .S(S[23]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1725 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_35), .S(S[22]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1721 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_36), .S(S[21]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1717 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_37), .S(S[20]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1713 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_38), .S(S[19]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1709 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_39), .S(S[18]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1705 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_40), .S(S[17]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1701 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_41), .S(S[16]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1697 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_42), .S(S[15]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1693 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_43), .S(S[14]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1689 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_44), .S(S[13]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1685 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_45), .S(S[12]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_1681 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_46), .S(S[11]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_1677 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(B[10]), .Cin(n_47), .S(S[10]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_1673 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), .B(), 
      .Cin(n_48), .S(S[9]), .P(), .G());
   Partial_Full_Adder__0_1669 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), .B(), 
      .Cin(n_49), .S(S[8]), .P(), .G());
   Partial_Full_Adder__0_1665 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_50), .S(S[7]), .P(), .G());
   Partial_Full_Adder__0_1661 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_51), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_1657 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_52), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_1653 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_53), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_1649 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_54), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_1645 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_55), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_1641 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_56), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_1637 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[26]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[9]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[8]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[7]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[6]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[5]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[4]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(A[3]), .A2(n_54), .ZN(n_53));
   AND2_X1 i_1_39 (.A1(A[2]), .A2(n_55), .ZN(n_54));
   AND2_X1 i_1_40 (.A1(A[1]), .A2(n_56), .ZN(n_55));
   AND2_X1 i_1_41 (.A1(Cin), .A2(A[0]), .ZN(n_56));
endmodule

module Partial_Full_Adder__0_1904(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1900(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1896(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1892(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1888(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1884(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1880(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1876(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1872(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1868(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1864(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1860(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1856(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1852(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1848(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1844(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_1840(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1836(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1832(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1828(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1824(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1820(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1816(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1812(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1808(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1804(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1800(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_1956(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_1904 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_32), .S(S[26]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_1900 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_33), .S(S[25]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_1896 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_34), .S(S[24]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_1892 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_35), .S(S[23]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_1888 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_36), .S(S[22]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_1884 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_37), .S(S[21]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_1880 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_38), .S(S[20]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_1876 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_39), .S(S[19]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_1872 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_40), .S(S[18]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_1868 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_41), .S(S[17]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_1864 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_42), .S(S[16]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_1860 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_43), .S(S[15]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_1856 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_44), .S(S[14]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_1852 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_45), .S(S[13]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_1848 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_46), .S(S[12]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_1844 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(B[11]), .Cin(n_47), .S(S[11]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_1840 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(), .Cin(n_48), .S(S[10]), .P(), .G());
   Partial_Full_Adder__0_1836 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), .B(), 
      .Cin(n_49), .S(S[9]), .P(), .G());
   Partial_Full_Adder__0_1832 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), .B(), 
      .Cin(n_50), .S(S[8]), .P(), .G());
   Partial_Full_Adder__0_1828 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_51), .S(S[7]), .P(), .G());
   Partial_Full_Adder__0_1824 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_52), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_1820 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_53), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_1816 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_54), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_1812 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_55), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_1808 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_56), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_1804 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_57), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_1800 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[27]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[10]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[9]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[8]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[7]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[6]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[5]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(A[4]), .A2(n_54), .ZN(n_53));
   AND2_X1 i_1_39 (.A1(A[3]), .A2(n_55), .ZN(n_54));
   AND2_X1 i_1_40 (.A1(A[2]), .A2(n_56), .ZN(n_55));
   AND2_X1 i_1_41 (.A1(A[1]), .A2(n_57), .ZN(n_56));
   AND2_X1 i_1_42 (.A1(Cin), .A2(A[0]), .ZN(n_57));
endmodule

module Partial_Full_Adder__0_2071(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2067(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2063(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2059(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2055(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2051(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2047(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2043(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2039(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2035(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2031(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2027(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2023(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2019(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2015(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2011(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2007(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2003(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1999(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1995(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1991(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1987(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1983(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1979(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1975(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1971(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1967(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_1963(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_2119(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_2071 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_32), .S(S[27]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2067 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_33), .S(S[26]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2063 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_34), .S(S[25]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2059 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_35), .S(S[24]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2055 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_36), .S(S[23]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2051 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_37), .S(S[22]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2047 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_38), .S(S[21]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2043 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_39), .S(S[20]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2039 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_40), .S(S[19]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2035 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_41), .S(S[18]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2031 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_42), .S(S[17]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2027 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_43), .S(S[16]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2023 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_44), .S(S[15]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2019 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_45), .S(S[14]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_2015 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_46), .S(S[13]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_2011 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(B[12]), .Cin(n_47), .S(S[12]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_2007 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(), .Cin(n_48), .S(S[11]), .P(), .G());
   Partial_Full_Adder__0_2003 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(), .Cin(n_49), .S(S[10]), .P(), .G());
   Partial_Full_Adder__0_1999 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), .B(), 
      .Cin(n_50), .S(S[9]), .P(), .G());
   Partial_Full_Adder__0_1995 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), .B(), 
      .Cin(n_51), .S(S[8]), .P(), .G());
   Partial_Full_Adder__0_1991 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_52), .S(S[7]), .P(), .G());
   Partial_Full_Adder__0_1987 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_53), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_1983 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_54), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_1979 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_55), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_1975 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_56), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_1971 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_57), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_1967 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_58), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_1963 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[28]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[11]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[10]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[9]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[8]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[7]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[6]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(A[5]), .A2(n_54), .ZN(n_53));
   AND2_X1 i_1_39 (.A1(A[4]), .A2(n_55), .ZN(n_54));
   AND2_X1 i_1_40 (.A1(A[3]), .A2(n_56), .ZN(n_55));
   AND2_X1 i_1_41 (.A1(A[2]), .A2(n_57), .ZN(n_56));
   AND2_X1 i_1_42 (.A1(A[1]), .A2(n_58), .ZN(n_57));
   AND2_X1 i_1_43 (.A1(Cin), .A2(A[0]), .ZN(n_58));
endmodule

module Partial_Full_Adder__0_2238(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2234(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2230(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2226(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2222(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2218(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2214(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2210(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2206(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2202(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2198(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2194(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2190(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2186(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2182(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2178(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2174(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2170(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2166(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2162(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2158(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2154(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2150(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2146(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2142(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2138(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2134(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2130(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2126(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_2282(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_2238 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_32), .S(S[28]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2234 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_33), .S(S[27]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2230 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2226 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_35), .S(S[25]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2222 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_36), .S(S[24]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2218 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_37), .S(S[23]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2214 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_38), .S(S[22]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2210 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_39), .S(S[21]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2206 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_40), .S(S[20]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2202 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_41), .S(S[19]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2198 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_42), .S(S[18]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2194 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_43), .S(S[17]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2190 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_44), .S(S[16]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2186 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_45), .S(S[15]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_2182 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_46), .S(S[14]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_2178 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(B[13]), .Cin(n_47), .S(S[13]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_2174 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(), .Cin(n_48), .S(S[12]), .P(), .G());
   Partial_Full_Adder__0_2170 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(), .Cin(n_49), .S(S[11]), .P(), .G());
   Partial_Full_Adder__0_2166 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(), .Cin(n_50), .S(S[10]), .P(), .G());
   Partial_Full_Adder__0_2162 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), .B(), 
      .Cin(n_51), .S(S[9]), .P(), .G());
   Partial_Full_Adder__0_2158 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), .B(), 
      .Cin(n_52), .S(S[8]), .P(), .G());
   Partial_Full_Adder__0_2154 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_53), .S(S[7]), .P(), .G());
   Partial_Full_Adder__0_2150 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_54), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_2146 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_55), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_2142 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_56), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_2138 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_57), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_2134 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_58), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_2130 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_59), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_2126 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[29]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[12]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[11]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[10]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[9]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[8]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[7]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(A[6]), .A2(n_54), .ZN(n_53));
   AND2_X1 i_1_39 (.A1(A[5]), .A2(n_55), .ZN(n_54));
   AND2_X1 i_1_40 (.A1(A[4]), .A2(n_56), .ZN(n_55));
   AND2_X1 i_1_41 (.A1(A[3]), .A2(n_57), .ZN(n_56));
   AND2_X1 i_1_42 (.A1(A[2]), .A2(n_58), .ZN(n_57));
   AND2_X1 i_1_43 (.A1(A[1]), .A2(n_59), .ZN(n_58));
   AND2_X1 i_1_44 (.A1(Cin), .A2(A[0]), .ZN(n_59));
endmodule

module Partial_Full_Adder__0_2405(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2401(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2397(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2393(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2389(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2385(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2381(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2377(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2373(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2369(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2365(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2361(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2357(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2353(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2349(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2345(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_2341(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2337(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2333(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2329(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2325(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2321(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2317(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2313(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2309(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2305(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2301(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2297(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2293(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_2289(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic__0_2445(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_15;

   Partial_Full_Adder__0_2405 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_32), .S(S[29]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_2401 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_33), .S(S[28]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_2397 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_34), .S(S[27]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_2393 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_35), .S(S[26]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_2389 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_36), .S(S[25]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_2385 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_37), .S(S[24]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_2381 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_38), .S(S[23]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_2377 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_39), .S(S[22]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_2373 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_40), .S(S[21]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_2369 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_41), .S(S[20]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_2365 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_42), .S(S[19]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_2361 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_43), .S(S[18]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_2357 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_44), .S(S[17]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_2353 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_45), .S(S[16]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_2349 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_46), .S(S[15]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_2345 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(B[14]), .Cin(n_47), .S(S[14]), .P(n_31), .G(n_30));
   Partial_Full_Adder__0_2341 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(), .Cin(n_48), .S(S[13]), .P(), .G());
   Partial_Full_Adder__0_2337 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(), .Cin(n_49), .S(S[12]), .P(), .G());
   Partial_Full_Adder__0_2333 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(), .Cin(n_50), .S(S[11]), .P(), .G());
   Partial_Full_Adder__0_2329 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(), .Cin(n_51), .S(S[10]), .P(), .G());
   Partial_Full_Adder__0_2325 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), .B(), 
      .Cin(n_52), .S(S[9]), .P(), .G());
   Partial_Full_Adder__0_2321 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), .B(), 
      .Cin(n_53), .S(S[8]), .P(), .G());
   Partial_Full_Adder__0_2317 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_54), .S(S[7]), .P(), .G());
   Partial_Full_Adder__0_2313 GEN_FULL_ADDERS_6_FULL_ADDER_INST (.A(A[6]), .B(), 
      .Cin(n_55), .S(S[6]), .P(), .G());
   Partial_Full_Adder__0_2309 GEN_FULL_ADDERS_5_FULL_ADDER_INST (.A(A[5]), .B(), 
      .Cin(n_56), .S(S[5]), .P(), .G());
   Partial_Full_Adder__0_2305 GEN_FULL_ADDERS_4_FULL_ADDER_INST (.A(A[4]), .B(), 
      .Cin(n_57), .S(S[4]), .P(), .G());
   Partial_Full_Adder__0_2301 GEN_FULL_ADDERS_3_FULL_ADDER_INST (.A(A[3]), .B(), 
      .Cin(n_58), .S(S[3]), .P(), .G());
   Partial_Full_Adder__0_2297 GEN_FULL_ADDERS_2_FULL_ADDER_INST (.A(A[2]), .B(), 
      .Cin(n_59), .S(S[2]), .P(), .G());
   Partial_Full_Adder__0_2293 GEN_FULL_ADDERS_1_FULL_ADDER_INST (.A(A[1]), .B(), 
      .Cin(n_60), .S(S[1]), .P(), .G());
   Partial_Full_Adder__0_2289 GEN_FULL_ADDERS_0_FULL_ADDER_INST (.A(A[0]), .B(), 
      .Cin(Cin), .S(S[0]), .P(), .G());
   OAI22_X1 i_0_0 (.A1(B[15]), .A2(n_0_1), .B1(n_0_0), .B2(S[15]), .ZN(overFlow));
   NAND2_X1 i_0_1 (.A1(A[15]), .A2(B[15]), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(S[15]), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(A[15]), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(S[30]));
   AOI21_X1 i_1_1 (.A(n_0), .B1(n_1), .B2(n_32), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(n_1_1), .ZN(n_32));
   AOI21_X1 i_1_3 (.A(n_2), .B1(n_3), .B2(n_33), .ZN(n_1_1));
   INV_X1 i_1_4 (.A(n_1_2), .ZN(n_33));
   AOI21_X1 i_1_5 (.A(n_4), .B1(n_5), .B2(n_34), .ZN(n_1_2));
   INV_X1 i_1_6 (.A(n_1_3), .ZN(n_34));
   AOI21_X1 i_1_7 (.A(n_6), .B1(n_7), .B2(n_35), .ZN(n_1_3));
   INV_X1 i_1_8 (.A(n_1_4), .ZN(n_35));
   AOI21_X1 i_1_9 (.A(n_8), .B1(n_9), .B2(n_36), .ZN(n_1_4));
   INV_X1 i_1_10 (.A(n_1_5), .ZN(n_36));
   AOI21_X1 i_1_11 (.A(n_10), .B1(n_11), .B2(n_37), .ZN(n_1_5));
   INV_X1 i_1_12 (.A(n_1_6), .ZN(n_37));
   AOI21_X1 i_1_13 (.A(n_12), .B1(n_13), .B2(n_38), .ZN(n_1_6));
   INV_X1 i_1_14 (.A(n_1_7), .ZN(n_38));
   AOI21_X1 i_1_15 (.A(n_14), .B1(n_15), .B2(n_39), .ZN(n_1_7));
   INV_X1 i_1_16 (.A(n_1_8), .ZN(n_39));
   AOI21_X1 i_1_17 (.A(n_16), .B1(n_17), .B2(n_40), .ZN(n_1_8));
   INV_X1 i_1_18 (.A(n_1_9), .ZN(n_40));
   AOI21_X1 i_1_19 (.A(n_18), .B1(n_19), .B2(n_41), .ZN(n_1_9));
   INV_X1 i_1_20 (.A(n_1_10), .ZN(n_41));
   AOI21_X1 i_1_21 (.A(n_20), .B1(n_21), .B2(n_42), .ZN(n_1_10));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_42));
   AOI21_X1 i_1_23 (.A(n_22), .B1(n_23), .B2(n_43), .ZN(n_1_11));
   INV_X1 i_1_24 (.A(n_1_12), .ZN(n_43));
   AOI21_X1 i_1_25 (.A(n_24), .B1(n_25), .B2(n_44), .ZN(n_1_12));
   INV_X1 i_1_26 (.A(n_1_13), .ZN(n_44));
   AOI21_X1 i_1_27 (.A(n_26), .B1(n_27), .B2(n_45), .ZN(n_1_13));
   INV_X1 i_1_28 (.A(n_1_14), .ZN(n_45));
   AOI21_X1 i_1_29 (.A(n_28), .B1(n_29), .B2(n_46), .ZN(n_1_14));
   INV_X1 i_1_30 (.A(n_1_15), .ZN(n_46));
   AOI21_X1 i_1_31 (.A(n_30), .B1(n_31), .B2(n_47), .ZN(n_1_15));
   AND2_X1 i_1_32 (.A1(A[13]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_1_33 (.A1(A[12]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_1_34 (.A1(A[11]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_1_35 (.A1(A[10]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_1_36 (.A1(A[9]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_1_37 (.A1(A[8]), .A2(n_53), .ZN(n_52));
   AND2_X1 i_1_38 (.A1(A[7]), .A2(n_54), .ZN(n_53));
   AND2_X1 i_1_39 (.A1(A[6]), .A2(n_55), .ZN(n_54));
   AND2_X1 i_1_40 (.A1(A[5]), .A2(n_56), .ZN(n_55));
   AND2_X1 i_1_41 (.A1(A[4]), .A2(n_57), .ZN(n_56));
   AND2_X1 i_1_42 (.A1(A[3]), .A2(n_58), .ZN(n_57));
   AND2_X1 i_1_43 (.A1(A[2]), .A2(n_59), .ZN(n_58));
   AND2_X1 i_1_44 (.A1(A[1]), .A2(n_60), .ZN(n_59));
   AND2_X1 i_1_45 (.A1(Cin), .A2(A[0]), .ZN(n_60));
endmodule

module Partial_Full_Adder__0_47(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_51(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_55(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_59(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_63(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_67(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_71(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_75(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_79(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_83(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_87(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_91(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_95(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_99(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_103(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_107(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_0_0 (.A(A), .B(B), .Z(P));
   XOR2_X1 i_0_1 (.A(P), .B(Cin), .Z(S));
   AND2_X1 i_0_2 (.A1(A), .A2(B), .ZN(G));
endmodule

module Partial_Full_Adder__0_111(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_115(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_119(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_123(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_127(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_131(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_135(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Partial_Full_Adder__0_139(A, B, Cin, S, P, G);
   input A;
   input B;
   input Cin;
   output S;
   output P;
   output G;

   XOR2_X1 i_1_0 (.A(A), .B(Cin), .Z(S));
endmodule

module Carry_Look_Ahead_generic(A, B, Cin, S, overFlow);
   input [31:0]A;
   input [31:0]B;
   input Cin;
   output [31:0]S;
   output overFlow;

   wire G;
   wire P;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;

   Partial_Full_Adder__0_47 GEN_FULL_ADDERS_30_FULL_ADDER_INST (.A(A[30]), 
      .B(B[30]), .Cin(n_30), .S(S[30]), .P(P), .G(G));
   Partial_Full_Adder__0_51 GEN_FULL_ADDERS_29_FULL_ADDER_INST (.A(A[29]), 
      .B(B[29]), .Cin(n_31), .S(S[29]), .P(n_1), .G(n_0));
   Partial_Full_Adder__0_55 GEN_FULL_ADDERS_28_FULL_ADDER_INST (.A(A[28]), 
      .B(B[28]), .Cin(n_32), .S(S[28]), .P(n_3), .G(n_2));
   Partial_Full_Adder__0_59 GEN_FULL_ADDERS_27_FULL_ADDER_INST (.A(A[27]), 
      .B(B[27]), .Cin(n_33), .S(S[27]), .P(n_5), .G(n_4));
   Partial_Full_Adder__0_63 GEN_FULL_ADDERS_26_FULL_ADDER_INST (.A(A[26]), 
      .B(B[26]), .Cin(n_34), .S(S[26]), .P(n_7), .G(n_6));
   Partial_Full_Adder__0_67 GEN_FULL_ADDERS_25_FULL_ADDER_INST (.A(A[25]), 
      .B(B[25]), .Cin(n_35), .S(S[25]), .P(n_9), .G(n_8));
   Partial_Full_Adder__0_71 GEN_FULL_ADDERS_24_FULL_ADDER_INST (.A(A[24]), 
      .B(B[24]), .Cin(n_36), .S(S[24]), .P(n_11), .G(n_10));
   Partial_Full_Adder__0_75 GEN_FULL_ADDERS_23_FULL_ADDER_INST (.A(A[23]), 
      .B(B[23]), .Cin(n_37), .S(S[23]), .P(n_13), .G(n_12));
   Partial_Full_Adder__0_79 GEN_FULL_ADDERS_22_FULL_ADDER_INST (.A(A[22]), 
      .B(B[22]), .Cin(n_38), .S(S[22]), .P(n_15), .G(n_14));
   Partial_Full_Adder__0_83 GEN_FULL_ADDERS_21_FULL_ADDER_INST (.A(A[21]), 
      .B(B[21]), .Cin(n_39), .S(S[21]), .P(n_17), .G(n_16));
   Partial_Full_Adder__0_87 GEN_FULL_ADDERS_20_FULL_ADDER_INST (.A(A[20]), 
      .B(B[20]), .Cin(n_40), .S(S[20]), .P(n_19), .G(n_18));
   Partial_Full_Adder__0_91 GEN_FULL_ADDERS_19_FULL_ADDER_INST (.A(A[19]), 
      .B(B[19]), .Cin(n_41), .S(S[19]), .P(n_21), .G(n_20));
   Partial_Full_Adder__0_95 GEN_FULL_ADDERS_18_FULL_ADDER_INST (.A(A[18]), 
      .B(B[18]), .Cin(n_42), .S(S[18]), .P(n_23), .G(n_22));
   Partial_Full_Adder__0_99 GEN_FULL_ADDERS_17_FULL_ADDER_INST (.A(A[17]), 
      .B(B[17]), .Cin(n_43), .S(S[17]), .P(n_25), .G(n_24));
   Partial_Full_Adder__0_103 GEN_FULL_ADDERS_16_FULL_ADDER_INST (.A(A[16]), 
      .B(B[16]), .Cin(n_44), .S(S[16]), .P(n_27), .G(n_26));
   Partial_Full_Adder__0_107 GEN_FULL_ADDERS_15_FULL_ADDER_INST (.A(A[15]), 
      .B(B[15]), .Cin(n_45), .S(S[15]), .P(n_29), .G(n_28));
   Partial_Full_Adder__0_111 GEN_FULL_ADDERS_14_FULL_ADDER_INST (.A(A[14]), 
      .B(), .Cin(n_46), .S(S[14]), .P(), .G());
   Partial_Full_Adder__0_115 GEN_FULL_ADDERS_13_FULL_ADDER_INST (.A(A[13]), 
      .B(), .Cin(n_47), .S(S[13]), .P(), .G());
   Partial_Full_Adder__0_119 GEN_FULL_ADDERS_12_FULL_ADDER_INST (.A(A[12]), 
      .B(), .Cin(n_48), .S(S[12]), .P(), .G());
   Partial_Full_Adder__0_123 GEN_FULL_ADDERS_11_FULL_ADDER_INST (.A(A[11]), 
      .B(), .Cin(n_49), .S(S[11]), .P(), .G());
   Partial_Full_Adder__0_127 GEN_FULL_ADDERS_10_FULL_ADDER_INST (.A(A[10]), 
      .B(), .Cin(n_50), .S(S[10]), .P(), .G());
   Partial_Full_Adder__0_131 GEN_FULL_ADDERS_9_FULL_ADDER_INST (.A(A[9]), .B(), 
      .Cin(n_51), .S(S[9]), .P(), .G());
   Partial_Full_Adder__0_135 GEN_FULL_ADDERS_8_FULL_ADDER_INST (.A(A[8]), .B(), 
      .Cin(n_52), .S(S[8]), .P(), .G());
   Partial_Full_Adder__0_139 GEN_FULL_ADDERS_7_FULL_ADDER_INST (.A(A[7]), .B(), 
      .Cin(n_53), .S(S[7]), .P(), .G());
   INV_X1 i_0_0 (.A(n_0_0), .ZN(S[31]));
   AOI21_X1 i_0_1 (.A(G), .B1(P), .B2(n_30), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(n_30));
   AOI21_X1 i_0_3 (.A(n_0), .B1(n_1), .B2(n_31), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(n_31));
   AOI21_X1 i_0_5 (.A(n_2), .B1(n_3), .B2(n_32), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_32));
   AOI21_X1 i_0_7 (.A(n_4), .B1(n_5), .B2(n_33), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_33));
   AOI21_X1 i_0_9 (.A(n_6), .B1(n_7), .B2(n_34), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(n_34));
   AOI21_X1 i_0_11 (.A(n_8), .B1(n_9), .B2(n_35), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(n_35));
   AOI21_X1 i_0_13 (.A(n_10), .B1(n_11), .B2(n_36), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(n_36));
   AOI21_X1 i_0_15 (.A(n_12), .B1(n_13), .B2(n_37), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(n_37));
   AOI21_X1 i_0_17 (.A(n_14), .B1(n_15), .B2(n_38), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(n_38));
   AOI21_X1 i_0_19 (.A(n_16), .B1(n_17), .B2(n_39), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(n_39));
   AOI21_X1 i_0_21 (.A(n_18), .B1(n_19), .B2(n_40), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(n_40));
   AOI21_X1 i_0_23 (.A(n_20), .B1(n_21), .B2(n_41), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(n_41));
   AOI21_X1 i_0_25 (.A(n_22), .B1(n_23), .B2(n_42), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(n_42));
   AOI21_X1 i_0_27 (.A(n_24), .B1(n_25), .B2(n_43), .ZN(n_0_13));
   INV_X1 i_0_28 (.A(n_0_14), .ZN(n_43));
   AOI21_X1 i_0_29 (.A(n_26), .B1(n_27), .B2(n_44), .ZN(n_0_14));
   INV_X1 i_0_30 (.A(n_0_15), .ZN(n_44));
   AOI21_X1 i_0_31 (.A(n_28), .B1(n_29), .B2(n_45), .ZN(n_0_15));
   AND2_X1 i_0_32 (.A1(A[14]), .A2(n_46), .ZN(n_45));
   AND2_X1 i_0_33 (.A1(A[13]), .A2(n_47), .ZN(n_46));
   AND2_X1 i_0_34 (.A1(A[12]), .A2(n_48), .ZN(n_47));
   AND2_X1 i_0_35 (.A1(A[11]), .A2(n_49), .ZN(n_48));
   AND2_X1 i_0_36 (.A1(A[10]), .A2(n_50), .ZN(n_49));
   AND2_X1 i_0_37 (.A1(A[9]), .A2(n_51), .ZN(n_50));
   AND2_X1 i_0_38 (.A1(A[8]), .A2(n_52), .ZN(n_51));
   AND2_X1 i_0_39 (.A1(A[7]), .A2(n_53), .ZN(n_52));
   NOR2_X1 i_0_40 (.A1(n_0_17), .A2(n_0_16), .ZN(n_53));
   NAND4_X1 i_0_41 (.A1(Cin), .A2(A[0]), .A3(A[1]), .A4(A[2]), .ZN(n_0_16));
   NAND4_X1 i_0_42 (.A1(A[3]), .A2(A[4]), .A3(A[5]), .A4(A[6]), .ZN(n_0_17));
endmodule

module AddandShift(A, B, Y, overflow);
   input [15:0]A;
   input [15:0]B;
   output [15:0]Y;
   output overflow;

   wire c;
   wire [31:0]\F[0] ;
   wire [31:0]\Z[15] ;
   wire [31:0]\Z[14] ;
   wire [31:0]\Z[13] ;
   wire [31:0]\Z[12] ;
   wire [31:0]\Z[11] ;
   wire [31:0]\Z[10] ;
   wire [31:0]\Z[9] ;
   wire [31:0]\Z[8] ;
   wire [31:0]\Z[7] ;
   wire [31:0]\Z[6] ;
   wire [31:0]\Z[5] ;
   wire [31:0]\Z[4] ;
   wire [31:0]\Z[3] ;
   wire [31:0]\Z[2] ;
   wire [31:0]\Z[1] ;
   wire [31:0]\Z[0] ;
   wire n_0_2;
   wire [31:0]\F[1] ;
   wire n_0_3;
   wire [31:0]\F[2] ;
   wire n_0_4;
   wire [31:0]\F[3] ;
   wire n_0_5;
   wire [31:0]\F[4] ;
   wire n_0_6;
   wire [31:0]\F[5] ;
   wire n_0_7;
   wire [31:0]\F[6] ;
   wire n_0_8;
   wire [31:0]\F[7] ;
   wire n_0_9;
   wire [31:0]\F[8] ;
   wire n_0_10;
   wire [31:0]\F[9] ;
   wire n_0_11;
   wire [31:0]\F[10] ;
   wire n_0_12;
   wire [31:0]\F[11] ;
   wire n_0_13;
   wire [31:0]\F[12] ;
   wire n_0_14;
   wire [31:0]\F[13] ;
   wire n_0_0;
   wire n_0_1;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;

   Carry_Look_Ahead_generic__0_326 p0 (.A({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, 
      uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      \Z[0] [15], \Z[0] [14], \Z[0] [13], \Z[0] [12], \Z[0] [11], \Z[0] [10], 
      \Z[0] [9], \Z[0] [8], \Z[0] [7], \Z[0] [6], \Z[0] [5], \Z[0] [4], 
      \Z[0] [3], \Z[0] [2], \Z[0] [1], uc_16}), .B({uc_17, uc_18, uc_19, uc_20, 
      uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, 
      uc_31, \Z[1] [16], \Z[1] [15], \Z[1] [14], \Z[1] [13], \Z[1] [12], 
      \Z[1] [11], \Z[1] [10], \Z[1] [9], \Z[1] [8], \Z[1] [7], \Z[1] [6], 
      \Z[1] [5], \Z[1] [4], \Z[1] [3], \Z[1] [2], \Z[1] [1], uc_32}), .Cin(), 
      .S({uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, 
      uc_43, uc_44, uc_45, uc_46, \F[0] [17], \F[0] [16], \F[0] [15], \F[0] [14], 
      \F[0] [13], \F[0] [12], \F[0] [11], \F[0] [10], \F[0] [9], \F[0] [8], 
      \F[0] [7], \F[0] [6], \F[0] [5], \F[0] [4], \F[0] [3], \F[0] [2], 
      \F[0] [1], uc_47}), .overFlow(c));
   MuxCustom__0_2447 L_15_li (.A({uc_48, A[15], A[14], A[13], A[12], A[11], 
      A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], uc_49, 
      uc_50, uc_51, uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, 
      uc_60, uc_61, uc_62, uc_63}), .Y({uc_64, \Z[15] [30], \Z[15] [29], 
      \Z[15] [28], \Z[15] [27], \Z[15] [26], \Z[15] [25], \Z[15] [24], 
      \Z[15] [23], \Z[15] [22], \Z[15] [21], \Z[15] [20], \Z[15] [19], 
      \Z[15] [18], \Z[15] [17], \Z[15] [16], \Z[15] [15], uc_65, uc_66, uc_67, 
      uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, 
      uc_78, uc_79}), .selector(B[15]));
   MuxCustom__0_2449 L_14_li (.A({uc_80, uc_81, A[15], A[14], A[13], A[12], 
      A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], 
      uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, 
      uc_92, uc_93, uc_94, uc_95}), .Y({uc_96, uc_97, \Z[14] [29], \Z[14] [28], 
      \Z[14] [27], \Z[14] [26], \Z[14] [25], \Z[14] [24], \Z[14] [23], 
      \Z[14] [22], \Z[14] [21], \Z[14] [20], \Z[14] [19], \Z[14] [18], 
      \Z[14] [17], \Z[14] [16], \Z[14] [15], \Z[14] [14], uc_98, uc_99, uc_100, 
      uc_101, uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, 
      uc_110, uc_111}), .selector(B[14]));
   MuxCustom__0_2451 L_13_li (.A({uc_112, uc_113, uc_114, A[15], A[14], A[13], 
      A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], 
      A[0], uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, 
      uc_123, uc_124, uc_125, uc_126, uc_127}), .Y({uc_128, uc_129, uc_130, 
      \Z[13] [28], \Z[13] [27], \Z[13] [26], \Z[13] [25], \Z[13] [24], 
      \Z[13] [23], \Z[13] [22], \Z[13] [21], \Z[13] [20], \Z[13] [19], 
      \Z[13] [18], \Z[13] [17], \Z[13] [16], \Z[13] [15], \Z[13] [14], 
      \Z[13] [13], uc_131, uc_132, uc_133, uc_134, uc_135, uc_136, uc_137, 
      uc_138, uc_139, uc_140, uc_141, uc_142, uc_143}), .selector(B[13]));
   MuxCustom__0_2453 L_12_li (.A({uc_144, uc_145, uc_146, uc_147, A[15], A[14], 
      A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], 
      A[1], A[0], uc_148, uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, uc_155, 
      uc_156, uc_157, uc_158, uc_159}), .Y({uc_160, uc_161, uc_162, uc_163, 
      \Z[12] [27], \Z[12] [26], \Z[12] [25], \Z[12] [24], \Z[12] [23], 
      \Z[12] [22], \Z[12] [21], \Z[12] [20], \Z[12] [19], \Z[12] [18], 
      \Z[12] [17], \Z[12] [16], \Z[12] [15], \Z[12] [14], \Z[12] [13], 
      \Z[12] [12], uc_164, uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, 
      uc_171, uc_172, uc_173, uc_174, uc_175}), .selector(B[12]));
   MuxCustom__0_2455 L_11_li (.A({uc_176, uc_177, uc_178, uc_179, uc_180, A[15], 
      A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], 
      A[3], A[2], A[1], A[0], uc_181, uc_182, uc_183, uc_184, uc_185, uc_186, 
      uc_187, uc_188, uc_189, uc_190, uc_191}), .Y({uc_192, uc_193, uc_194, 
      uc_195, uc_196, \Z[11] [26], \Z[11] [25], \Z[11] [24], \Z[11] [23], 
      \Z[11] [22], \Z[11] [21], \Z[11] [20], \Z[11] [19], \Z[11] [18], 
      \Z[11] [17], \Z[11] [16], \Z[11] [15], \Z[11] [14], \Z[11] [13], 
      \Z[11] [12], \Z[11] [11], uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, 
      uc_203, uc_204, uc_205, uc_206, uc_207}), .selector(B[11]));
   MuxCustom__0_2457 L_10_li (.A({uc_208, uc_209, uc_210, uc_211, uc_212, uc_213, 
      A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], 
      A[4], A[3], A[2], A[1], A[0], uc_214, uc_215, uc_216, uc_217, uc_218, 
      uc_219, uc_220, uc_221, uc_222, uc_223}), .Y({uc_224, uc_225, uc_226, 
      uc_227, uc_228, uc_229, \Z[10] [25], \Z[10] [24], \Z[10] [23], \Z[10] [22], 
      \Z[10] [21], \Z[10] [20], \Z[10] [19], \Z[10] [18], \Z[10] [17], 
      \Z[10] [16], \Z[10] [15], \Z[10] [14], \Z[10] [13], \Z[10] [12], 
      \Z[10] [11], \Z[10] [10], uc_230, uc_231, uc_232, uc_233, uc_234, uc_235, 
      uc_236, uc_237, uc_238, uc_239}), .selector(B[10]));
   MuxCustom__0_2459 L_9_li (.A({uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, 
      uc_246, A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], 
      A[5], A[4], A[3], A[2], A[1], A[0], uc_247, uc_248, uc_249, uc_250, uc_251, 
      uc_252, uc_253, uc_254, uc_255}), .Y({uc_256, uc_257, uc_258, uc_259, 
      uc_260, uc_261, uc_262, \Z[9] [24], \Z[9] [23], \Z[9] [22], \Z[9] [21], 
      \Z[9] [20], \Z[9] [19], \Z[9] [18], \Z[9] [17], \Z[9] [16], \Z[9] [15], 
      \Z[9] [14], \Z[9] [13], \Z[9] [12], \Z[9] [11], \Z[9] [10], \Z[9] [9], 
      uc_263, uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271}), 
      .selector(B[9]));
   MuxCustom__0_2461 L_8_li (.A({uc_272, uc_273, uc_274, uc_275, uc_276, uc_277, 
      uc_278, uc_279, A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], 
      A[6], A[5], A[4], A[3], A[2], A[1], A[0], uc_280, uc_281, uc_282, uc_283, 
      uc_284, uc_285, uc_286, uc_287}), .Y({uc_288, uc_289, uc_290, uc_291, 
      uc_292, uc_293, uc_294, uc_295, \Z[8] [23], \Z[8] [22], \Z[8] [21], 
      \Z[8] [20], \Z[8] [19], \Z[8] [18], \Z[8] [17], \Z[8] [16], \Z[8] [15], 
      \Z[8] [14], \Z[8] [13], \Z[8] [12], \Z[8] [11], \Z[8] [10], \Z[8] [9], 
      \Z[8] [8], uc_296, uc_297, uc_298, uc_299, uc_300, uc_301, uc_302, uc_303}), 
      .selector(B[8]));
   MuxCustom__0_2463 L_7_li (.A({uc_304, uc_305, uc_306, uc_307, uc_308, uc_309, 
      uc_310, uc_311, uc_312, A[15], A[14], A[13], A[12], A[11], A[10], A[9], 
      A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], uc_313, uc_314, 
      uc_315, uc_316, uc_317, uc_318, uc_319}), .Y({uc_320, uc_321, uc_322, 
      uc_323, uc_324, uc_325, uc_326, uc_327, uc_328, \Z[7] [22], \Z[7] [21], 
      \Z[7] [20], \Z[7] [19], \Z[7] [18], \Z[7] [17], \Z[7] [16], \Z[7] [15], 
      \Z[7] [14], \Z[7] [13], \Z[7] [12], \Z[7] [11], \Z[7] [10], \Z[7] [9], 
      \Z[7] [8], \Z[7] [7], uc_329, uc_330, uc_331, uc_332, uc_333, uc_334, 
      uc_335}), .selector(B[7]));
   MuxCustom__0_2465 L_6_li (.A({uc_336, uc_337, uc_338, uc_339, uc_340, uc_341, 
      uc_342, uc_343, uc_344, uc_345, A[15], A[14], A[13], A[12], A[11], A[10], 
      A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], uc_346, uc_347, 
      uc_348, uc_349, uc_350, uc_351}), .Y({uc_352, uc_353, uc_354, uc_355, 
      uc_356, uc_357, uc_358, uc_359, uc_360, uc_361, \Z[6] [21], \Z[6] [20], 
      \Z[6] [19], \Z[6] [18], \Z[6] [17], \Z[6] [16], \Z[6] [15], \Z[6] [14], 
      \Z[6] [13], \Z[6] [12], \Z[6] [11], \Z[6] [10], \Z[6] [9], \Z[6] [8], 
      \Z[6] [7], \Z[6] [6], uc_362, uc_363, uc_364, uc_365, uc_366, uc_367}), 
      .selector(B[6]));
   MuxCustom__0_2467 L_5_li (.A({uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, 
      uc_374, uc_375, uc_376, uc_377, uc_378, A[15], A[14], A[13], A[12], A[11], 
      A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], uc_379, 
      uc_380, uc_381, uc_382, uc_383}), .Y({uc_384, uc_385, uc_386, uc_387, 
      uc_388, uc_389, uc_390, uc_391, uc_392, uc_393, uc_394, \Z[5] [20], 
      \Z[5] [19], \Z[5] [18], \Z[5] [17], \Z[5] [16], \Z[5] [15], \Z[5] [14], 
      \Z[5] [13], \Z[5] [12], \Z[5] [11], \Z[5] [10], \Z[5] [9], \Z[5] [8], 
      \Z[5] [7], \Z[5] [6], \Z[5] [5], uc_395, uc_396, uc_397, uc_398, uc_399}), 
      .selector(B[5]));
   MuxCustom__0_2469 L_4_li (.A({uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, 
      uc_406, uc_407, uc_408, uc_409, uc_410, uc_411, A[15], A[14], A[13], A[12], 
      A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0], 
      uc_412, uc_413, uc_414, uc_415}), .Y({uc_416, uc_417, uc_418, uc_419, 
      uc_420, uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, \Z[4] [19], 
      \Z[4] [18], \Z[4] [17], \Z[4] [16], \Z[4] [15], \Z[4] [14], \Z[4] [13], 
      \Z[4] [12], \Z[4] [11], \Z[4] [10], \Z[4] [9], \Z[4] [8], \Z[4] [7], 
      \Z[4] [6], \Z[4] [5], \Z[4] [4], uc_428, uc_429, uc_430, uc_431}), 
      .selector(B[4]));
   MuxCustom__0_2471 L_3_li (.A({uc_432, uc_433, uc_434, uc_435, uc_436, uc_437, 
      uc_438, uc_439, uc_440, uc_441, uc_442, uc_443, uc_444, A[15], A[14], 
      A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], 
      A[1], A[0], uc_445, uc_446, uc_447}), .Y({uc_448, uc_449, uc_450, uc_451, 
      uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, uc_459, uc_460, 
      \Z[3] [18], \Z[3] [17], \Z[3] [16], \Z[3] [15], \Z[3] [14], \Z[3] [13], 
      \Z[3] [12], \Z[3] [11], \Z[3] [10], \Z[3] [9], \Z[3] [8], \Z[3] [7], 
      \Z[3] [6], \Z[3] [5], \Z[3] [4], \Z[3] [3], uc_461, uc_462, uc_463}), 
      .selector(B[3]));
   MuxCustom__0_2473 L_2_li (.A({uc_464, uc_465, uc_466, uc_467, uc_468, uc_469, 
      uc_470, uc_471, uc_472, uc_473, uc_474, uc_475, uc_476, uc_477, A[15], 
      A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], A[4], 
      A[3], A[2], A[1], A[0], uc_478, uc_479}), .Y({uc_480, uc_481, uc_482, 
      uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489, uc_490, uc_491, 
      uc_492, uc_493, \Z[2] [17], \Z[2] [16], \Z[2] [15], \Z[2] [14], \Z[2] [13], 
      \Z[2] [12], \Z[2] [11], \Z[2] [10], \Z[2] [9], \Z[2] [8], \Z[2] [7], 
      \Z[2] [6], \Z[2] [5], \Z[2] [4], \Z[2] [3], \Z[2] [2], uc_494, uc_495}), 
      .selector(B[2]));
   MuxCustom__0_2475 L_1_li (.A({uc_496, uc_497, uc_498, uc_499, uc_500, uc_501, 
      uc_502, uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, uc_509, uc_510, 
      A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], 
      A[4], A[3], A[2], A[1], A[0], uc_511}), .Y({uc_512, uc_513, uc_514, uc_515, 
      uc_516, uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524, 
      uc_525, uc_526, \Z[1] [16], \Z[1] [15], \Z[1] [14], \Z[1] [13], \Z[1] [12], 
      \Z[1] [11], \Z[1] [10], \Z[1] [9], \Z[1] [8], \Z[1] [7], \Z[1] [6], 
      \Z[1] [5], \Z[1] [4], \Z[1] [3], \Z[1] [2], \Z[1] [1], uc_527}), .selector(
      B[1]));
   MuxCustom L_0_li (.A({uc_528, uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, 
      uc_535, uc_536, uc_537, uc_538, uc_539, uc_540, uc_541, uc_542, uc_543, 
      A[15], A[14], A[13], A[12], A[11], A[10], A[9], A[8], A[7], A[6], A[5], 
      A[4], A[3], A[2], A[1], A[0]}), .Y({uc_544, uc_545, uc_546, uc_547, uc_548, 
      uc_549, uc_550, uc_551, uc_552, uc_553, uc_554, uc_555, uc_556, uc_557, 
      uc_558, uc_559, \Z[0] [15], \Z[0] [14], \Z[0] [13], \Z[0] [12], \Z[0] [11], 
      \Z[0] [10], \Z[0] [9], \Z[0] [8], \Z[0] [7], \Z[0] [6], \Z[0] [5], 
      \Z[0] [4], \Z[0] [3], \Z[0] [2], \Z[0] [1], \Z[0] [0]}), .selector(B[0]));
   Carry_Look_Ahead_generic__0_489 p_0_pi (.A({uc_560, uc_561, uc_562, uc_563, 
      uc_564, uc_565, uc_566, uc_567, uc_568, uc_569, uc_570, uc_571, uc_572, 
      uc_573, \F[0] [17], \F[0] [16], \F[0] [15], \F[0] [14], \F[0] [13], 
      \F[0] [12], \F[0] [11], \F[0] [10], \F[0] [9], \F[0] [8], \F[0] [7], 
      \F[0] [6], \F[0] [5], \F[0] [4], \F[0] [3], \F[0] [2], \F[0] [1], 
      \Z[0] [0]}), .B({uc_574, uc_575, uc_576, uc_577, uc_578, uc_579, uc_580, 
      uc_581, uc_582, uc_583, uc_584, uc_585, uc_586, uc_587, \Z[2] [17], 
      \Z[2] [16], \Z[2] [15], \Z[2] [14], \Z[2] [13], \Z[2] [12], \Z[2] [11], 
      \Z[2] [10], \Z[2] [9], \Z[2] [8], \Z[2] [7], \Z[2] [6], \Z[2] [5], 
      \Z[2] [4], \Z[2] [3], \Z[2] [2], uc_588, uc_589}), .Cin(c), .S({uc_590, 
      uc_591, uc_592, uc_593, uc_594, uc_595, uc_596, uc_597, uc_598, uc_599, 
      uc_600, uc_601, uc_602, \F[1] [18], \F[1] [17], \F[1] [16], \F[1] [15], 
      \F[1] [14], \F[1] [13], \F[1] [12], \F[1] [11], \F[1] [10], \F[1] [9], 
      \F[1] [8], \F[1] [7], \F[1] [6], \F[1] [5], \F[1] [4], \F[1] [3], 
      \F[1] [2], \F[1] [1], \F[1] [0]}), .overFlow(n_0_2));
   Carry_Look_Ahead_generic__0_652 p_1_pi (.A({uc_603, uc_604, uc_605, uc_606, 
      uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, uc_615, 
      \F[1] [18], \F[1] [17], \F[1] [16], \F[1] [15], \F[1] [14], \F[1] [13], 
      \F[1] [12], \F[1] [11], \F[1] [10], \F[1] [9], \F[1] [8], \F[1] [7], 
      \F[1] [6], \F[1] [5], \F[1] [4], \F[1] [3], \F[1] [2], \F[1] [1], 
      \F[1] [0]}), .B({uc_616, uc_617, uc_618, uc_619, uc_620, uc_621, uc_622, 
      uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, \Z[3] [18], \Z[3] [17], 
      \Z[3] [16], \Z[3] [15], \Z[3] [14], \Z[3] [13], \Z[3] [12], \Z[3] [11], 
      \Z[3] [10], \Z[3] [9], \Z[3] [8], \Z[3] [7], \Z[3] [6], \Z[3] [5], 
      \Z[3] [4], \Z[3] [3], uc_629, uc_630, uc_631}), .Cin(n_0_2), .S({uc_632, 
      uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, uc_639, uc_640, uc_641, 
      uc_642, uc_643, \F[2] [19], \F[2] [18], \F[2] [17], \F[2] [16], \F[2] [15], 
      \F[2] [14], \F[2] [13], \F[2] [12], \F[2] [11], \F[2] [10], \F[2] [9], 
      \F[2] [8], \F[2] [7], \F[2] [6], \F[2] [5], \F[2] [4], \F[2] [3], 
      \F[2] [2], \F[2] [1], \F[2] [0]}), .overFlow(n_0_3));
   Carry_Look_Ahead_generic__0_815 p_2_pi (.A({uc_644, uc_645, uc_646, uc_647, 
      uc_648, uc_649, uc_650, uc_651, uc_652, uc_653, uc_654, uc_655, \F[2] [19], 
      \F[2] [18], \F[2] [17], \F[2] [16], \F[2] [15], \F[2] [14], \F[2] [13], 
      \F[2] [12], \F[2] [11], \F[2] [10], \F[2] [9], \F[2] [8], \F[2] [7], 
      \F[2] [6], \F[2] [5], \F[2] [4], \F[2] [3], \F[2] [2], \F[2] [1], 
      \F[2] [0]}), .B({uc_656, uc_657, uc_658, uc_659, uc_660, uc_661, uc_662, 
      uc_663, uc_664, uc_665, uc_666, uc_667, \Z[4] [19], \Z[4] [18], \Z[4] [17], 
      \Z[4] [16], \Z[4] [15], \Z[4] [14], \Z[4] [13], \Z[4] [12], \Z[4] [11], 
      \Z[4] [10], \Z[4] [9], \Z[4] [8], \Z[4] [7], \Z[4] [6], \Z[4] [5], 
      \Z[4] [4], uc_668, uc_669, uc_670, uc_671}), .Cin(n_0_3), .S({uc_672, 
      uc_673, uc_674, uc_675, uc_676, uc_677, uc_678, uc_679, uc_680, uc_681, 
      uc_682, \F[3] [20], \F[3] [19], \F[3] [18], \F[3] [17], \F[3] [16], 
      \F[3] [15], \F[3] [14], \F[3] [13], \F[3] [12], \F[3] [11], \F[3] [10], 
      \F[3] [9], \F[3] [8], \F[3] [7], \F[3] [6], \F[3] [5], \F[3] [4], 
      \F[3] [3], \F[3] [2], \F[3] [1], \F[3] [0]}), .overFlow(n_0_4));
   Carry_Look_Ahead_generic__0_978 p_3_pi (.A({uc_683, uc_684, uc_685, uc_686, 
      uc_687, uc_688, uc_689, uc_690, uc_691, uc_692, uc_693, \F[3] [20], 
      \F[3] [19], \F[3] [18], \F[3] [17], \F[3] [16], \F[3] [15], \F[3] [14], 
      \F[3] [13], \F[3] [12], \F[3] [11], \F[3] [10], \F[3] [9], \F[3] [8], 
      \F[3] [7], \F[3] [6], \F[3] [5], \F[3] [4], \F[3] [3], \F[3] [2], 
      \F[3] [1], \F[3] [0]}), .B({uc_694, uc_695, uc_696, uc_697, uc_698, uc_699, 
      uc_700, uc_701, uc_702, uc_703, uc_704, \Z[5] [20], \Z[5] [19], \Z[5] [18], 
      \Z[5] [17], \Z[5] [16], \Z[5] [15], \Z[5] [14], \Z[5] [13], \Z[5] [12], 
      \Z[5] [11], \Z[5] [10], \Z[5] [9], \Z[5] [8], \Z[5] [7], \Z[5] [6], 
      \Z[5] [5], uc_705, uc_706, uc_707, uc_708, uc_709}), .Cin(n_0_4), .S({
      uc_710, uc_711, uc_712, uc_713, uc_714, uc_715, uc_716, uc_717, uc_718, 
      uc_719, \F[4] [21], \F[4] [20], \F[4] [19], \F[4] [18], \F[4] [17], 
      \F[4] [16], \F[4] [15], \F[4] [14], \F[4] [13], \F[4] [12], \F[4] [11], 
      \F[4] [10], \F[4] [9], \F[4] [8], \F[4] [7], \F[4] [6], \F[4] [5], 
      \F[4] [4], \F[4] [3], \F[4] [2], \F[4] [1], \F[4] [0]}), .overFlow(n_0_5));
   Carry_Look_Ahead_generic__0_1141 p_4_pi (.A({uc_720, uc_721, uc_722, uc_723, 
      uc_724, uc_725, uc_726, uc_727, uc_728, uc_729, \F[4] [21], \F[4] [20], 
      \F[4] [19], \F[4] [18], \F[4] [17], \F[4] [16], \F[4] [15], \F[4] [14], 
      \F[4] [13], \F[4] [12], \F[4] [11], \F[4] [10], \F[4] [9], \F[4] [8], 
      \F[4] [7], \F[4] [6], \F[4] [5], \F[4] [4], \F[4] [3], \F[4] [2], 
      \F[4] [1], \F[4] [0]}), .B({uc_730, uc_731, uc_732, uc_733, uc_734, uc_735, 
      uc_736, uc_737, uc_738, uc_739, \Z[6] [21], \Z[6] [20], \Z[6] [19], 
      \Z[6] [18], \Z[6] [17], \Z[6] [16], \Z[6] [15], \Z[6] [14], \Z[6] [13], 
      \Z[6] [12], \Z[6] [11], \Z[6] [10], \Z[6] [9], \Z[6] [8], \Z[6] [7], 
      \Z[6] [6], uc_740, uc_741, uc_742, uc_743, uc_744, uc_745}), .Cin(n_0_5), 
      .S({uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752, uc_753, uc_754, 
      \F[5] [22], \F[5] [21], \F[5] [20], \F[5] [19], \F[5] [18], \F[5] [17], 
      \F[5] [16], \F[5] [15], \F[5] [14], \F[5] [13], \F[5] [12], \F[5] [11], 
      \F[5] [10], \F[5] [9], \F[5] [8], \F[5] [7], \F[5] [6], \F[5] [5], 
      \F[5] [4], \F[5] [3], \F[5] [2], \F[5] [1], \F[5] [0]}), .overFlow(n_0_6));
   Carry_Look_Ahead_generic__0_1304 p_5_pi (.A({uc_755, uc_756, uc_757, uc_758, 
      uc_759, uc_760, uc_761, uc_762, uc_763, \F[5] [22], \F[5] [21], \F[5] [20], 
      \F[5] [19], \F[5] [18], \F[5] [17], \F[5] [16], \F[5] [15], \F[5] [14], 
      \F[5] [13], \F[5] [12], \F[5] [11], \F[5] [10], \F[5] [9], \F[5] [8], 
      \F[5] [7], \F[5] [6], \F[5] [5], \F[5] [4], \F[5] [3], \F[5] [2], 
      \F[5] [1], \F[5] [0]}), .B({uc_764, uc_765, uc_766, uc_767, uc_768, uc_769, 
      uc_770, uc_771, uc_772, \Z[7] [22], \Z[7] [21], \Z[7] [20], \Z[7] [19], 
      \Z[7] [18], \Z[7] [17], \Z[7] [16], \Z[7] [15], \Z[7] [14], \Z[7] [13], 
      \Z[7] [12], \Z[7] [11], \Z[7] [10], \Z[7] [9], \Z[7] [8], \Z[7] [7], 
      uc_773, uc_774, uc_775, uc_776, uc_777, uc_778, uc_779}), .Cin(n_0_6), 
      .S({uc_780, uc_781, uc_782, uc_783, uc_784, uc_785, uc_786, uc_787, 
      \F[6] [23], \F[6] [22], \F[6] [21], \F[6] [20], \F[6] [19], \F[6] [18], 
      \F[6] [17], \F[6] [16], \F[6] [15], \F[6] [14], \F[6] [13], \F[6] [12], 
      \F[6] [11], \F[6] [10], \F[6] [9], \F[6] [8], \F[6] [7], \F[6] [6], 
      \F[6] [5], \F[6] [4], \F[6] [3], \F[6] [2], \F[6] [1], \F[6] [0]}), 
      .overFlow(n_0_7));
   Carry_Look_Ahead_generic__0_1467 p_6_pi (.A({uc_788, uc_789, uc_790, uc_791, 
      uc_792, uc_793, uc_794, uc_795, \F[6] [23], \F[6] [22], \F[6] [21], 
      \F[6] [20], \F[6] [19], \F[6] [18], \F[6] [17], \F[6] [16], \F[6] [15], 
      \F[6] [14], \F[6] [13], \F[6] [12], \F[6] [11], \F[6] [10], \F[6] [9], 
      \F[6] [8], \F[6] [7], \F[6] [6], \F[6] [5], \F[6] [4], \F[6] [3], 
      \F[6] [2], \F[6] [1], \F[6] [0]}), .B({uc_796, uc_797, uc_798, uc_799, 
      uc_800, uc_801, uc_802, uc_803, \Z[8] [23], \Z[8] [22], \Z[8] [21], 
      \Z[8] [20], \Z[8] [19], \Z[8] [18], \Z[8] [17], \Z[8] [16], \Z[8] [15], 
      \Z[8] [14], \Z[8] [13], \Z[8] [12], \Z[8] [11], \Z[8] [10], \Z[8] [9], 
      \Z[8] [8], uc_804, uc_805, uc_806, uc_807, uc_808, uc_809, uc_810, uc_811}), 
      .Cin(n_0_7), .S({uc_812, uc_813, uc_814, uc_815, uc_816, uc_817, uc_818, 
      \F[7] [24], \F[7] [23], \F[7] [22], \F[7] [21], \F[7] [20], \F[7] [19], 
      \F[7] [18], \F[7] [17], \F[7] [16], \F[7] [15], \F[7] [14], \F[7] [13], 
      \F[7] [12], \F[7] [11], \F[7] [10], \F[7] [9], \F[7] [8], \F[7] [7], 
      \F[7] [6], \F[7] [5], \F[7] [4], \F[7] [3], \F[7] [2], \F[7] [1], 
      \F[7] [0]}), .overFlow(n_0_8));
   Carry_Look_Ahead_generic__0_1630 p_7_pi (.A({uc_819, uc_820, uc_821, uc_822, 
      uc_823, uc_824, uc_825, \F[7] [24], \F[7] [23], \F[7] [22], \F[7] [21], 
      \F[7] [20], \F[7] [19], \F[7] [18], \F[7] [17], \F[7] [16], \F[7] [15], 
      \F[7] [14], \F[7] [13], \F[7] [12], \F[7] [11], \F[7] [10], \F[7] [9], 
      \F[7] [8], \F[7] [7], \F[7] [6], \F[7] [5], \F[7] [4], \F[7] [3], 
      \F[7] [2], \F[7] [1], \F[7] [0]}), .B({uc_826, uc_827, uc_828, uc_829, 
      uc_830, uc_831, uc_832, \Z[9] [24], \Z[9] [23], \Z[9] [22], \Z[9] [21], 
      \Z[9] [20], \Z[9] [19], \Z[9] [18], \Z[9] [17], \Z[9] [16], \Z[9] [15], 
      \Z[9] [14], \Z[9] [13], \Z[9] [12], \Z[9] [11], \Z[9] [10], \Z[9] [9], 
      uc_833, uc_834, uc_835, uc_836, uc_837, uc_838, uc_839, uc_840, uc_841}), 
      .Cin(n_0_8), .S({uc_842, uc_843, uc_844, uc_845, uc_846, uc_847, 
      \F[8] [25], \F[8] [24], \F[8] [23], \F[8] [22], \F[8] [21], \F[8] [20], 
      \F[8] [19], \F[8] [18], \F[8] [17], \F[8] [16], \F[8] [15], \F[8] [14], 
      \F[8] [13], \F[8] [12], \F[8] [11], \F[8] [10], \F[8] [9], \F[8] [8], 
      \F[8] [7], \F[8] [6], \F[8] [5], \F[8] [4], \F[8] [3], \F[8] [2], 
      \F[8] [1], \F[8] [0]}), .overFlow(n_0_9));
   Carry_Look_Ahead_generic__0_1793 p_8_pi (.A({uc_848, uc_849, uc_850, uc_851, 
      uc_852, uc_853, \F[8] [25], \F[8] [24], \F[8] [23], \F[8] [22], \F[8] [21], 
      \F[8] [20], \F[8] [19], \F[8] [18], \F[8] [17], \F[8] [16], \F[8] [15], 
      \F[8] [14], \F[8] [13], \F[8] [12], \F[8] [11], \F[8] [10], \F[8] [9], 
      \F[8] [8], \F[8] [7], \F[8] [6], \F[8] [5], \F[8] [4], \F[8] [3], 
      \F[8] [2], \F[8] [1], \F[8] [0]}), .B({uc_854, uc_855, uc_856, uc_857, 
      uc_858, uc_859, \Z[10] [25], \Z[10] [24], \Z[10] [23], \Z[10] [22], 
      \Z[10] [21], \Z[10] [20], \Z[10] [19], \Z[10] [18], \Z[10] [17], 
      \Z[10] [16], \Z[10] [15], \Z[10] [14], \Z[10] [13], \Z[10] [12], 
      \Z[10] [11], \Z[10] [10], uc_860, uc_861, uc_862, uc_863, uc_864, uc_865, 
      uc_866, uc_867, uc_868, uc_869}), .Cin(n_0_9), .S({uc_870, uc_871, uc_872, 
      uc_873, uc_874, \F[9] [26], \F[9] [25], \F[9] [24], \F[9] [23], \F[9] [22], 
      \F[9] [21], \F[9] [20], \F[9] [19], \F[9] [18], \F[9] [17], \F[9] [16], 
      \F[9] [15], \F[9] [14], \F[9] [13], \F[9] [12], \F[9] [11], \F[9] [10], 
      \F[9] [9], \F[9] [8], \F[9] [7], \F[9] [6], \F[9] [5], \F[9] [4], 
      \F[9] [3], \F[9] [2], \F[9] [1], \F[9] [0]}), .overFlow(n_0_10));
   Carry_Look_Ahead_generic__0_1956 p_9_pi (.A({uc_875, uc_876, uc_877, uc_878, 
      uc_879, \F[9] [26], \F[9] [25], \F[9] [24], \F[9] [23], \F[9] [22], 
      \F[9] [21], \F[9] [20], \F[9] [19], \F[9] [18], \F[9] [17], \F[9] [16], 
      \F[9] [15], \F[9] [14], \F[9] [13], \F[9] [12], \F[9] [11], \F[9] [10], 
      \F[9] [9], \F[9] [8], \F[9] [7], \F[9] [6], \F[9] [5], \F[9] [4], 
      \F[9] [3], \F[9] [2], \F[9] [1], \F[9] [0]}), .B({uc_880, uc_881, uc_882, 
      uc_883, uc_884, \Z[11] [26], \Z[11] [25], \Z[11] [24], \Z[11] [23], 
      \Z[11] [22], \Z[11] [21], \Z[11] [20], \Z[11] [19], \Z[11] [18], 
      \Z[11] [17], \Z[11] [16], \Z[11] [15], \Z[11] [14], \Z[11] [13], 
      \Z[11] [12], \Z[11] [11], uc_885, uc_886, uc_887, uc_888, uc_889, uc_890, 
      uc_891, uc_892, uc_893, uc_894, uc_895}), .Cin(n_0_10), .S({uc_896, uc_897, 
      uc_898, uc_899, \F[10] [27], \F[10] [26], \F[10] [25], \F[10] [24], 
      \F[10] [23], \F[10] [22], \F[10] [21], \F[10] [20], \F[10] [19], 
      \F[10] [18], \F[10] [17], \F[10] [16], \F[10] [15], \F[10] [14], 
      \F[10] [13], \F[10] [12], \F[10] [11], \F[10] [10], \F[10] [9], \F[10] [8], 
      \F[10] [7], \F[10] [6], \F[10] [5], \F[10] [4], \F[10] [3], \F[10] [2], 
      \F[10] [1], \F[10] [0]}), .overFlow(n_0_11));
   Carry_Look_Ahead_generic__0_2119 p_10_pi (.A({uc_900, uc_901, uc_902, uc_903, 
      \F[10] [27], \F[10] [26], \F[10] [25], \F[10] [24], \F[10] [23], 
      \F[10] [22], \F[10] [21], \F[10] [20], \F[10] [19], \F[10] [18], 
      \F[10] [17], \F[10] [16], \F[10] [15], \F[10] [14], \F[10] [13], 
      \F[10] [12], \F[10] [11], \F[10] [10], \F[10] [9], \F[10] [8], \F[10] [7], 
      \F[10] [6], \F[10] [5], \F[10] [4], \F[10] [3], \F[10] [2], \F[10] [1], 
      \F[10] [0]}), .B({uc_904, uc_905, uc_906, uc_907, \Z[12] [27], \Z[12] [26], 
      \Z[12] [25], \Z[12] [24], \Z[12] [23], \Z[12] [22], \Z[12] [21], 
      \Z[12] [20], \Z[12] [19], \Z[12] [18], \Z[12] [17], \Z[12] [16], 
      \Z[12] [15], \Z[12] [14], \Z[12] [13], \Z[12] [12], uc_908, uc_909, uc_910, 
      uc_911, uc_912, uc_913, uc_914, uc_915, uc_916, uc_917, uc_918, uc_919}), 
      .Cin(n_0_11), .S({uc_920, uc_921, uc_922, \F[11] [28], \F[11] [27], 
      \F[11] [26], \F[11] [25], \F[11] [24], \F[11] [23], \F[11] [22], 
      \F[11] [21], \F[11] [20], \F[11] [19], \F[11] [18], \F[11] [17], 
      \F[11] [16], \F[11] [15], \F[11] [14], \F[11] [13], \F[11] [12], 
      \F[11] [11], \F[11] [10], \F[11] [9], \F[11] [8], \F[11] [7], \F[11] [6], 
      \F[11] [5], \F[11] [4], \F[11] [3], \F[11] [2], \F[11] [1], \F[11] [0]}), 
      .overFlow(n_0_12));
   Carry_Look_Ahead_generic__0_2282 p_11_pi (.A({uc_923, uc_924, uc_925, 
      \F[11] [28], \F[11] [27], \F[11] [26], \F[11] [25], \F[11] [24], 
      \F[11] [23], \F[11] [22], \F[11] [21], \F[11] [20], \F[11] [19], 
      \F[11] [18], \F[11] [17], \F[11] [16], \F[11] [15], \F[11] [14], 
      \F[11] [13], \F[11] [12], \F[11] [11], \F[11] [10], \F[11] [9], \F[11] [8], 
      \F[11] [7], \F[11] [6], \F[11] [5], \F[11] [4], \F[11] [3], \F[11] [2], 
      \F[11] [1], \F[11] [0]}), .B({uc_926, uc_927, uc_928, \Z[13] [28], 
      \Z[13] [27], \Z[13] [26], \Z[13] [25], \Z[13] [24], \Z[13] [23], 
      \Z[13] [22], \Z[13] [21], \Z[13] [20], \Z[13] [19], \Z[13] [18], 
      \Z[13] [17], \Z[13] [16], \Z[13] [15], \Z[13] [14], \Z[13] [13], uc_929, 
      uc_930, uc_931, uc_932, uc_933, uc_934, uc_935, uc_936, uc_937, uc_938, 
      uc_939, uc_940, uc_941}), .Cin(n_0_12), .S({uc_942, uc_943, \F[12] [29], 
      \F[12] [28], \F[12] [27], \F[12] [26], \F[12] [25], \F[12] [24], 
      \F[12] [23], \F[12] [22], \F[12] [21], \F[12] [20], \F[12] [19], 
      \F[12] [18], \F[12] [17], \F[12] [16], \F[12] [15], \F[12] [14], 
      \F[12] [13], \F[12] [12], \F[12] [11], \F[12] [10], \F[12] [9], \F[12] [8], 
      \F[12] [7], \F[12] [6], \F[12] [5], \F[12] [4], \F[12] [3], \F[12] [2], 
      \F[12] [1], \F[12] [0]}), .overFlow(n_0_13));
   Carry_Look_Ahead_generic__0_2445 p_12_pi (.A({uc_944, uc_945, \F[12] [29], 
      \F[12] [28], \F[12] [27], \F[12] [26], \F[12] [25], \F[12] [24], 
      \F[12] [23], \F[12] [22], \F[12] [21], \F[12] [20], \F[12] [19], 
      \F[12] [18], \F[12] [17], \F[12] [16], \F[12] [15], \F[12] [14], 
      \F[12] [13], \F[12] [12], \F[12] [11], \F[12] [10], \F[12] [9], \F[12] [8], 
      \F[12] [7], \F[12] [6], \F[12] [5], \F[12] [4], \F[12] [3], \F[12] [2], 
      \F[12] [1], \F[12] [0]}), .B({uc_946, uc_947, \Z[14] [29], \Z[14] [28], 
      \Z[14] [27], \Z[14] [26], \Z[14] [25], \Z[14] [24], \Z[14] [23], 
      \Z[14] [22], \Z[14] [21], \Z[14] [20], \Z[14] [19], \Z[14] [18], 
      \Z[14] [17], \Z[14] [16], \Z[14] [15], \Z[14] [14], uc_948, uc_949, uc_950, 
      uc_951, uc_952, uc_953, uc_954, uc_955, uc_956, uc_957, uc_958, uc_959, 
      uc_960, uc_961}), .Cin(n_0_13), .S({uc_962, \F[13] [30], \F[13] [29], 
      \F[13] [28], \F[13] [27], \F[13] [26], \F[13] [25], \F[13] [24], 
      \F[13] [23], \F[13] [22], \F[13] [21], \F[13] [20], \F[13] [19], 
      \F[13] [18], \F[13] [17], \F[13] [16], \F[13] [15], \F[13] [14], 
      \F[13] [13], \F[13] [12], \F[13] [11], \F[13] [10], \F[13] [9], \F[13] [8], 
      \F[13] [7], \F[13] [6], \F[13] [5], \F[13] [4], \F[13] [3], \F[13] [2], 
      \F[13] [1], \F[13] [0]}), .overFlow(n_0_14));
   Carry_Look_Ahead_generic p_13_pi (.A({uc_963, \F[13] [30], \F[13] [29], 
      \F[13] [28], \F[13] [27], \F[13] [26], \F[13] [25], \F[13] [24], 
      \F[13] [23], \F[13] [22], \F[13] [21], \F[13] [20], \F[13] [19], 
      \F[13] [18], \F[13] [17], \F[13] [16], \F[13] [15], \F[13] [14], 
      \F[13] [13], \F[13] [12], \F[13] [11], \F[13] [10], \F[13] [9], \F[13] [8], 
      \F[13] [7], \F[13] [6], \F[13] [5], \F[13] [4], \F[13] [3], \F[13] [2], 
      \F[13] [1], \F[13] [0]}), .B({uc_964, \Z[15] [30], \Z[15] [29], 
      \Z[15] [28], \Z[15] [27], \Z[15] [26], \Z[15] [25], \Z[15] [24], 
      \Z[15] [23], \Z[15] [22], \Z[15] [21], \Z[15] [20], \Z[15] [19], 
      \Z[15] [18], \Z[15] [17], \Z[15] [16], \Z[15] [15], uc_965, uc_966, uc_967, 
      uc_968, uc_969, uc_970, uc_971, uc_972, uc_973, uc_974, uc_975, uc_976, 
      uc_977, uc_978, uc_979}), .Cin(n_0_14), .S({n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, n_0_1, n_0_0, Y[15], Y[14], Y[13], Y[12], Y[11], 
      Y[10], Y[9], Y[8], Y[7], Y[6], Y[5], Y[4], Y[3], Y[2], Y[1], Y[0], uc_980, 
      uc_981, uc_982, uc_983, uc_984, uc_985, uc_986}), .overFlow());
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(overflow));
   OAI33_X1 i_0_0_1 (.A1(n_0_0_4), .A2(n_0_0_2), .A3(n_0_0_5), .B1(n_0_0_3), 
      .B2(n_0_0_1), .B3(n_0_21), .ZN(n_0_0_0));
   OR4_X1 i_0_0_2 (.A1(n_0_19), .A2(n_0_18), .A3(n_0_20), .A4(n_0_17), .ZN(
      n_0_0_1));
   NAND4_X1 i_0_0_3 (.A1(n_0_19), .A2(n_0_18), .A3(n_0_20), .A4(n_0_17), 
      .ZN(n_0_0_2));
   OR4_X1 i_0_0_4 (.A1(n_0_16), .A2(n_0_15), .A3(n_0_1), .A4(n_0_0), .ZN(n_0_0_3));
   NAND4_X1 i_0_0_5 (.A1(n_0_16), .A2(n_0_15), .A3(n_0_1), .A4(n_0_0), .ZN(
      n_0_0_4));
   INV_X1 i_0_0_6 (.A(n_0_21), .ZN(n_0_0_5));
endmodule
