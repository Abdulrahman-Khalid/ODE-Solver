/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 12:51:44 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3743315520 */

module datapath(addr_T, p_0);
   input [31:0]addr_T;
   output [31:0]p_0;

   HA_X1 i_1 (.A(addr_T[1]), .B(addr_T[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_2 (.A(addr_T[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_3 (.A(addr_T[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_4 (.A(addr_T[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_5 (.A(addr_T[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_6 (.A(addr_T[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_7 (.A(addr_T[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_8 (.A(addr_T[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_9 (.A(addr_T[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_10 (.A(addr_T[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(addr_T[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(addr_T[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(addr_T[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(addr_T[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(addr_T[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(addr_T[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(addr_T[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(addr_T[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(addr_T[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_20 (.A(addr_T[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_21 (.A(addr_T[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_22 (.A(addr_T[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_23 (.A(addr_T[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_24 (.A(addr_T[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_25 (.A(addr_T[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_26 (.A(addr_T[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_27 (.A(addr_T[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_28 (.A(addr_T[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_29 (.A(addr_T[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_30 (.A(addr_T[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_0 (.A(addr_T[31]), .B(n_29), .Z(p_0[31]));
   INV_X1 i_31 (.A(addr_T[0]), .ZN(p_0[0]));
endmodule

module datapath__0_144(addr_output, p_0);
   input [31:0]addr_output;
   output [31:0]p_0;

   HA_X1 i_0 (.A(addr_output[1]), .B(addr_output[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_1 (.A(addr_output[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_2 (.A(addr_output[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_3 (.A(addr_output[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_4 (.A(addr_output[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_5 (.A(addr_output[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_6 (.A(addr_output[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_7 (.A(addr_output[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_8 (.A(addr_output[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_9 (.A(addr_output[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(addr_output[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(addr_output[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(addr_output[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(addr_output[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(addr_output[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(addr_output[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(addr_output[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(addr_output[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(addr_output[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_10 (.A(addr_output[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_20 (.A(addr_output[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_21 (.A(addr_output[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_22 (.A(addr_output[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_23 (.A(addr_output[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_24 (.A(addr_output[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_25 (.A(addr_output[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_26 (.A(addr_output[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_27 (.A(addr_output[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_28 (.A(addr_output[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_29 (.A(addr_output[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_30 (.A(addr_output[31]), .B(n_29), .Z(p_0[31]));
   INV_X1 i_31 (.A(addr_output[0]), .ZN(p_0[0]));
endmodule

module IO_Output(enable_output_IO, CLK, RST, end_T_address, end_Output_address, 
      memory_data, CPU_Bus, memory_address, done_output_data);
   input enable_output_IO;
   input CLK;
   input RST;
   input [31:0]end_T_address;
   input [31:0]end_Output_address;
   input [63:0]memory_data;
   output [31:0]CPU_Bus;
   output [31:0]memory_address;
   output done_output_data;

   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire [1:0]state_reg;
   wire n_0_269;
   wire n_0_270;
   wire n_0_272;
   wire n_0_274;
   wire n_0_276;
   wire n_0_278;
   wire n_0_280;
   wire n_0_282;
   wire n_0_284;
   wire n_0_286;
   wire n_0_288;
   wire n_0_290;
   wire n_0_292;
   wire n_0_294;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire [1:0]state;
   wire n_0_119;
   wire n_0_232;
   wire n_0_0_0;
   wire n_0_231;
   wire n_0_0_1;
   wire n_0_230;
   wire n_0_0_2;
   wire n_0_229;
   wire n_0_0_3;
   wire n_0_228;
   wire n_0_0_4;
   wire n_0_227;
   wire n_0_0_5;
   wire n_0_226;
   wire n_0_0_6;
   wire n_0_225;
   wire n_0_0_7;
   wire n_0_224;
   wire n_0_0_8;
   wire n_0_223;
   wire n_0_0_9;
   wire n_0_222;
   wire n_0_0_10;
   wire n_0_221;
   wire n_0_0_11;
   wire n_0_220;
   wire n_0_0_12;
   wire n_0_219;
   wire n_0_0_13;
   wire n_0_218;
   wire n_0_0_14;
   wire n_0_217;
   wire n_0_0_15;
   wire n_0_216;
   wire n_0_0_16;
   wire n_0_215;
   wire n_0_0_17;
   wire n_0_214;
   wire n_0_0_18;
   wire n_0_213;
   wire n_0_0_19;
   wire n_0_212;
   wire n_0_0_20;
   wire n_0_211;
   wire n_0_0_21;
   wire n_0_210;
   wire n_0_0_22;
   wire n_0_209;
   wire n_0_0_23;
   wire n_0_208;
   wire n_0_0_24;
   wire n_0_207;
   wire n_0_0_25;
   wire n_0_206;
   wire n_0_0_26;
   wire n_0_205;
   wire n_0_0_27;
   wire n_0_204;
   wire n_0_0_28;
   wire n_0_203;
   wire n_0_0_29;
   wire n_0_202;
   wire n_0_0_30;
   wire n_0_200;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_117;
   wire n_0_0_35;
   wire n_0_198;
   wire n_0_197;
   wire n_0_196;
   wire n_0_195;
   wire n_0_194;
   wire n_0_193;
   wire n_0_192;
   wire n_0_191;
   wire n_0_190;
   wire n_0_189;
   wire n_0_188;
   wire n_0_187;
   wire n_0_186;
   wire n_0_185;
   wire n_0_184;
   wire n_0_183;
   wire n_0_182;
   wire n_0_181;
   wire n_0_180;
   wire n_0_179;
   wire n_0_178;
   wire n_0_177;
   wire n_0_176;
   wire n_0_175;
   wire n_0_174;
   wire n_0_173;
   wire n_0_172;
   wire n_0_171;
   wire n_0_170;
   wire n_0_169;
   wire n_0_168;
   wire n_0_167;
   wire n_0_0_36;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_199;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire eq;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_249;
   wire n_0_0_87;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_0_88;
   wire n_0_254;
   wire n_0_0_89;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_0_90;
   wire n_0_258;
   wire n_0_0_91;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_0_92;
   wire n_0_262;
   wire n_0_0_93;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_0_94;
   wire n_0_266;
   wire n_0_0_95;
   wire n_0_267;
   wire n_0_268;
   wire n_0_271;
   wire n_0_0_96;
   wire n_0_273;
   wire n_0_0_97;
   wire n_0_275;
   wire n_0_277;
   wire n_0_279;
   wire n_0_0_98;
   wire n_0_281;
   wire n_0_0_99;
   wire n_0_283;
   wire n_0_285;
   wire n_0_287;
   wire n_0_0_100;
   wire n_0_289;
   wire n_0_0_101;
   wire n_0_291;
   wire n_0_0_102;
   wire n_0_293;
   wire n_0_118;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_295;
   wire n_0_201;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;

   DFFR_X1 done_output_data_reg (.D(state_reg[1]), .RN(n_0_295), .CK(n_0_201), 
      .Q(done_output_data), .QN());
   CLKGATETST_X1 clk_gate_memory_address_reg (.CK(CLK), .E(eq), .SE(1'b0), 
      .GCK(n_0_3));
   DFF_X1 \memory_address_reg[31]  (.D(n_0_293), .CK(n_0_3), .Q(
      memory_address[31]), .QN());
   DFF_X1 \memory_address_reg[30]  (.D(n_0_291), .CK(n_0_3), .Q(
      memory_address[30]), .QN());
   DFF_X1 \memory_address_reg[29]  (.D(n_0_289), .CK(n_0_3), .Q(
      memory_address[29]), .QN());
   DFF_X1 \memory_address_reg[28]  (.D(n_0_287), .CK(n_0_3), .Q(
      memory_address[28]), .QN());
   DFF_X1 \memory_address_reg[27]  (.D(n_0_285), .CK(n_0_3), .Q(
      memory_address[27]), .QN());
   DFF_X1 \memory_address_reg[26]  (.D(n_0_283), .CK(n_0_3), .Q(
      memory_address[26]), .QN());
   DFF_X1 \memory_address_reg[25]  (.D(n_0_281), .CK(n_0_3), .Q(
      memory_address[25]), .QN());
   DFF_X1 \memory_address_reg[24]  (.D(n_0_279), .CK(n_0_3), .Q(
      memory_address[24]), .QN());
   DFF_X1 \memory_address_reg[23]  (.D(n_0_277), .CK(n_0_3), .Q(
      memory_address[23]), .QN());
   DFF_X1 \memory_address_reg[22]  (.D(n_0_275), .CK(n_0_3), .Q(
      memory_address[22]), .QN());
   DFF_X1 \memory_address_reg[21]  (.D(n_0_273), .CK(n_0_3), .Q(
      memory_address[21]), .QN());
   DFF_X1 \memory_address_reg[20]  (.D(n_0_271), .CK(n_0_3), .Q(
      memory_address[20]), .QN());
   DFF_X1 \memory_address_reg[19]  (.D(n_0_268), .CK(n_0_3), .Q(
      memory_address[19]), .QN());
   DFF_X1 \memory_address_reg[18]  (.D(n_0_267), .CK(n_0_3), .Q(
      memory_address[18]), .QN());
   DFF_X1 \memory_address_reg[17]  (.D(n_0_266), .CK(n_0_3), .Q(
      memory_address[17]), .QN());
   DFF_X1 \memory_address_reg[16]  (.D(n_0_265), .CK(n_0_3), .Q(
      memory_address[16]), .QN());
   DFF_X1 \memory_address_reg[15]  (.D(n_0_264), .CK(n_0_3), .Q(
      memory_address[15]), .QN());
   DFF_X1 \memory_address_reg[14]  (.D(n_0_263), .CK(n_0_3), .Q(
      memory_address[14]), .QN());
   DFF_X1 \memory_address_reg[13]  (.D(n_0_262), .CK(n_0_3), .Q(
      memory_address[13]), .QN());
   DFF_X1 \memory_address_reg[12]  (.D(n_0_261), .CK(n_0_3), .Q(
      memory_address[12]), .QN());
   DFF_X1 \memory_address_reg[11]  (.D(n_0_260), .CK(n_0_3), .Q(
      memory_address[11]), .QN());
   DFF_X1 \memory_address_reg[10]  (.D(n_0_259), .CK(n_0_3), .Q(
      memory_address[10]), .QN());
   DFF_X1 \memory_address_reg[9]  (.D(n_0_258), .CK(n_0_3), .Q(memory_address[9]), 
      .QN());
   DFF_X1 \memory_address_reg[8]  (.D(n_0_257), .CK(n_0_3), .Q(memory_address[8]), 
      .QN());
   DFF_X1 \memory_address_reg[7]  (.D(n_0_256), .CK(n_0_3), .Q(memory_address[7]), 
      .QN());
   DFF_X1 \memory_address_reg[6]  (.D(n_0_255), .CK(n_0_3), .Q(memory_address[6]), 
      .QN());
   DFF_X1 \memory_address_reg[5]  (.D(n_0_254), .CK(n_0_3), .Q(memory_address[5]), 
      .QN());
   DFF_X1 \memory_address_reg[4]  (.D(n_0_253), .CK(n_0_3), .Q(memory_address[4]), 
      .QN());
   DFF_X1 \memory_address_reg[3]  (.D(n_0_252), .CK(n_0_3), .Q(memory_address[3]), 
      .QN());
   DFF_X1 \memory_address_reg[2]  (.D(n_0_251), .CK(n_0_3), .Q(memory_address[2]), 
      .QN());
   DFF_X1 \memory_address_reg[1]  (.D(n_0_250), .CK(n_0_3), .Q(memory_address[1]), 
      .QN());
   DFF_X1 \memory_address_reg[0]  (.D(n_0_249), .CK(n_0_3), .Q(memory_address[0]), 
      .QN());
   datapath i_0_3 (.addr_T({n_0_85, n_0_86, n_0_87, n_0_88, n_0_89, n_0_90, 
      n_0_91, n_0_92, n_0_93, n_0_94, n_0_95, n_0_96, n_0_97, n_0_98, n_0_99, 
      n_0_100, n_0_101, n_0_102, n_0_103, n_0_104, n_0_105, n_0_106, n_0_107, 
      n_0_108, n_0_109, n_0_110, n_0_111, n_0_112, n_0_113, n_0_114, n_0_115, 
      n_0_116}), .p_0({n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, 
      n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, 
      n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
      n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4}));
   DFFRS_X1 \memory_address_reg[31]__0  (.D(n_0_167), .RN(n_0_248), .SN(n_0_166), 
      .CK(n_0_201), .Q(memory_address[31]), .QN());
   DFFRS_X1 \memory_address_reg[30]__0  (.D(n_0_168), .RN(n_0_247), .SN(n_0_165), 
      .CK(n_0_201), .Q(memory_address[30]), .QN());
   DFFRS_X1 \memory_address_reg[29]__0  (.D(n_0_169), .RN(n_0_246), .SN(n_0_164), 
      .CK(n_0_201), .Q(memory_address[29]), .QN());
   DFFRS_X1 \memory_address_reg[28]__0  (.D(n_0_170), .RN(n_0_245), .SN(n_0_163), 
      .CK(n_0_201), .Q(memory_address[28]), .QN());
   DFFRS_X1 \memory_address_reg[27]__0  (.D(n_0_171), .RN(n_0_244), .SN(n_0_162), 
      .CK(n_0_201), .Q(memory_address[27]), .QN());
   DFFRS_X1 \memory_address_reg[26]__0  (.D(n_0_172), .RN(n_0_243), .SN(n_0_161), 
      .CK(n_0_201), .Q(memory_address[26]), .QN());
   DFFRS_X1 \memory_address_reg[25]__0  (.D(n_0_173), .RN(n_0_242), .SN(n_0_160), 
      .CK(n_0_201), .Q(memory_address[25]), .QN());
   DFFRS_X1 \memory_address_reg[24]__0  (.D(n_0_174), .RN(n_0_241), .SN(n_0_159), 
      .CK(n_0_201), .Q(memory_address[24]), .QN());
   DFFRS_X1 \memory_address_reg[23]__0  (.D(n_0_175), .RN(n_0_240), .SN(n_0_158), 
      .CK(n_0_201), .Q(memory_address[23]), .QN());
   DFFRS_X1 \memory_address_reg[22]__0  (.D(n_0_176), .RN(n_0_239), .SN(n_0_157), 
      .CK(n_0_201), .Q(memory_address[22]), .QN());
   DFFRS_X1 \memory_address_reg[21]__0  (.D(n_0_177), .RN(n_0_238), .SN(n_0_156), 
      .CK(n_0_201), .Q(memory_address[21]), .QN());
   DFFRS_X1 \memory_address_reg[20]__0  (.D(n_0_178), .RN(n_0_237), .SN(n_0_155), 
      .CK(n_0_201), .Q(memory_address[20]), .QN());
   DFFRS_X1 \memory_address_reg[19]__0  (.D(n_0_179), .RN(n_0_236), .SN(n_0_154), 
      .CK(n_0_201), .Q(memory_address[19]), .QN());
   DFFRS_X1 \memory_address_reg[18]__0  (.D(n_0_180), .RN(n_0_235), .SN(n_0_153), 
      .CK(n_0_201), .Q(memory_address[18]), .QN());
   DFFRS_X1 \memory_address_reg[17]__0  (.D(n_0_181), .RN(n_0_234), .SN(n_0_152), 
      .CK(n_0_201), .Q(memory_address[17]), .QN());
   DFFRS_X1 \memory_address_reg[16]__0  (.D(n_0_182), .RN(n_0_233), .SN(n_0_151), 
      .CK(n_0_201), .Q(memory_address[16]), .QN());
   DFFRS_X1 \memory_address_reg[15]__0  (.D(n_0_183), .RN(n_0_199), .SN(n_0_150), 
      .CK(n_0_201), .Q(memory_address[15]), .QN());
   DFFRS_X1 \memory_address_reg[14]__0  (.D(n_0_184), .RN(n_0_134), .SN(n_0_149), 
      .CK(n_0_201), .Q(memory_address[14]), .QN());
   DFFRS_X1 \memory_address_reg[13]__0  (.D(n_0_185), .RN(n_0_133), .SN(n_0_148), 
      .CK(n_0_201), .Q(memory_address[13]), .QN());
   DFFRS_X1 \memory_address_reg[12]__0  (.D(n_0_186), .RN(n_0_132), .SN(n_0_147), 
      .CK(n_0_201), .Q(memory_address[12]), .QN());
   DFFRS_X1 \memory_address_reg[11]__0  (.D(n_0_187), .RN(n_0_131), .SN(n_0_146), 
      .CK(n_0_201), .Q(memory_address[11]), .QN());
   DFFRS_X1 \memory_address_reg[10]__0  (.D(n_0_188), .RN(n_0_130), .SN(n_0_145), 
      .CK(n_0_201), .Q(memory_address[10]), .QN());
   DFFRS_X1 \memory_address_reg[9]__0  (.D(n_0_189), .RN(n_0_129), .SN(n_0_144), 
      .CK(n_0_201), .Q(memory_address[9]), .QN());
   DFFRS_X1 \memory_address_reg[8]__0  (.D(n_0_190), .RN(n_0_128), .SN(n_0_143), 
      .CK(n_0_201), .Q(memory_address[8]), .QN());
   DFFRS_X1 \memory_address_reg[7]__0  (.D(n_0_191), .RN(n_0_127), .SN(n_0_142), 
      .CK(n_0_201), .Q(memory_address[7]), .QN());
   DFFRS_X1 \memory_address_reg[6]__0  (.D(n_0_192), .RN(n_0_126), .SN(n_0_141), 
      .CK(n_0_201), .Q(memory_address[6]), .QN());
   DFFRS_X1 \memory_address_reg[5]__0  (.D(n_0_193), .RN(n_0_125), .SN(n_0_140), 
      .CK(n_0_201), .Q(memory_address[5]), .QN());
   DFFRS_X1 \memory_address_reg[4]__0  (.D(n_0_194), .RN(n_0_124), .SN(n_0_139), 
      .CK(n_0_201), .Q(memory_address[4]), .QN());
   DFFRS_X1 \memory_address_reg[3]__0  (.D(n_0_195), .RN(n_0_123), .SN(n_0_138), 
      .CK(n_0_201), .Q(memory_address[3]), .QN());
   DFFRS_X1 \memory_address_reg[2]__0  (.D(n_0_196), .RN(n_0_122), .SN(n_0_137), 
      .CK(n_0_201), .Q(memory_address[2]), .QN());
   DFFRS_X1 \memory_address_reg[1]__0  (.D(n_0_197), .RN(n_0_121), .SN(n_0_136), 
      .CK(n_0_201), .Q(memory_address[1]), .QN());
   DFFRS_X1 \memory_address_reg[0]__0  (.D(n_0_198), .RN(n_0_120), .SN(n_0_135), 
      .CK(n_0_201), .Q(memory_address[0]), .QN());
   DFF_X1 \CPU_Bus_reg[31]  (.D(n_0_200), .CK(n_0_201), .Q(CPU_Bus[31]), .QN());
   DFF_X1 \CPU_Bus_reg[30]  (.D(n_0_202), .CK(n_0_201), .Q(CPU_Bus[30]), .QN());
   DFF_X1 \CPU_Bus_reg[29]  (.D(n_0_203), .CK(n_0_201), .Q(CPU_Bus[29]), .QN());
   DFF_X1 \CPU_Bus_reg[28]  (.D(n_0_204), .CK(n_0_201), .Q(CPU_Bus[28]), .QN());
   DFF_X1 \CPU_Bus_reg[27]  (.D(n_0_205), .CK(n_0_201), .Q(CPU_Bus[27]), .QN());
   DFF_X1 \CPU_Bus_reg[26]  (.D(n_0_206), .CK(n_0_201), .Q(CPU_Bus[26]), .QN());
   DFF_X1 \CPU_Bus_reg[25]  (.D(n_0_207), .CK(n_0_201), .Q(CPU_Bus[25]), .QN());
   DFF_X1 \CPU_Bus_reg[24]  (.D(n_0_208), .CK(n_0_201), .Q(CPU_Bus[24]), .QN());
   DFF_X1 \CPU_Bus_reg[23]  (.D(n_0_209), .CK(n_0_201), .Q(CPU_Bus[23]), .QN());
   DFF_X1 \CPU_Bus_reg[22]  (.D(n_0_210), .CK(n_0_201), .Q(CPU_Bus[22]), .QN());
   DFF_X1 \CPU_Bus_reg[21]  (.D(n_0_211), .CK(n_0_201), .Q(CPU_Bus[21]), .QN());
   DFF_X1 \CPU_Bus_reg[20]  (.D(n_0_212), .CK(n_0_201), .Q(CPU_Bus[20]), .QN());
   DFF_X1 \CPU_Bus_reg[19]  (.D(n_0_213), .CK(n_0_201), .Q(CPU_Bus[19]), .QN());
   DFF_X1 \CPU_Bus_reg[18]  (.D(n_0_214), .CK(n_0_201), .Q(CPU_Bus[18]), .QN());
   DFF_X1 \CPU_Bus_reg[17]  (.D(n_0_215), .CK(n_0_201), .Q(CPU_Bus[17]), .QN());
   DFF_X1 \CPU_Bus_reg[16]  (.D(n_0_216), .CK(n_0_201), .Q(CPU_Bus[16]), .QN());
   DFF_X1 \CPU_Bus_reg[15]  (.D(n_0_217), .CK(n_0_201), .Q(CPU_Bus[15]), .QN());
   DFF_X1 \CPU_Bus_reg[14]  (.D(n_0_218), .CK(n_0_201), .Q(CPU_Bus[14]), .QN());
   DFF_X1 \CPU_Bus_reg[13]  (.D(n_0_219), .CK(n_0_201), .Q(CPU_Bus[13]), .QN());
   DFF_X1 \CPU_Bus_reg[12]  (.D(n_0_220), .CK(n_0_201), .Q(CPU_Bus[12]), .QN());
   DFF_X1 \CPU_Bus_reg[11]  (.D(n_0_221), .CK(n_0_201), .Q(CPU_Bus[11]), .QN());
   DFF_X1 \CPU_Bus_reg[10]  (.D(n_0_222), .CK(n_0_201), .Q(CPU_Bus[10]), .QN());
   DFF_X1 \CPU_Bus_reg[9]  (.D(n_0_223), .CK(n_0_201), .Q(CPU_Bus[9]), .QN());
   DFF_X1 \CPU_Bus_reg[8]  (.D(n_0_224), .CK(n_0_201), .Q(CPU_Bus[8]), .QN());
   DFF_X1 \CPU_Bus_reg[7]  (.D(n_0_225), .CK(n_0_201), .Q(CPU_Bus[7]), .QN());
   DFF_X1 \CPU_Bus_reg[6]  (.D(n_0_226), .CK(n_0_201), .Q(CPU_Bus[6]), .QN());
   DFF_X1 \CPU_Bus_reg[5]  (.D(n_0_227), .CK(n_0_201), .Q(CPU_Bus[5]), .QN());
   DFF_X1 \CPU_Bus_reg[4]  (.D(n_0_228), .CK(n_0_201), .Q(CPU_Bus[4]), .QN());
   DFF_X1 \CPU_Bus_reg[3]  (.D(n_0_229), .CK(n_0_201), .Q(CPU_Bus[3]), .QN());
   DFF_X1 \CPU_Bus_reg[2]  (.D(n_0_230), .CK(n_0_201), .Q(CPU_Bus[2]), .QN());
   DFF_X1 \CPU_Bus_reg[1]  (.D(n_0_231), .CK(n_0_201), .Q(CPU_Bus[1]), .QN());
   DFF_X1 \CPU_Bus_reg[0]  (.D(n_0_232), .CK(n_0_201), .Q(CPU_Bus[0]), .QN());
   DFF_X1 \state_reg[1]  (.D(done_output_data), .CK(CLK), .Q(state_reg[1]), 
      .QN());
   DFF_X1 \state_reg[0]  (.D(state[0]), .CK(CLK), .Q(state_reg[0]), .QN());
   CLKGATETST_X1 clk_gate_addr_output_reg (.CK(CLK), .E(n_0_119), .SE(1'b0), 
      .GCK(n_0_269));
   DFFR_X1 \addr_output_reg[31]  (.D(n_0_83), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_270), .QN());
   DFFR_X1 \addr_output_reg[30]  (.D(n_0_82), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_272), .QN());
   DFFR_X1 \addr_output_reg[29]  (.D(n_0_81), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_274), .QN());
   DFFR_X1 \addr_output_reg[28]  (.D(n_0_80), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_276), .QN());
   DFFR_X1 \addr_output_reg[27]  (.D(n_0_79), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_278), .QN());
   DFFR_X1 \addr_output_reg[26]  (.D(n_0_78), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_280), .QN());
   DFFR_X1 \addr_output_reg[25]  (.D(n_0_77), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_282), .QN());
   DFFR_X1 \addr_output_reg[24]  (.D(n_0_76), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_284), .QN());
   DFFR_X1 \addr_output_reg[23]  (.D(n_0_75), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_286), .QN());
   DFFR_X1 \addr_output_reg[22]  (.D(n_0_74), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_288), .QN());
   DFFR_X1 \addr_output_reg[21]  (.D(n_0_73), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_290), .QN());
   DFFR_X1 \addr_output_reg[20]  (.D(n_0_72), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_292), .QN());
   DFFR_X1 \addr_output_reg[19]  (.D(n_0_71), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_294), .QN());
   DFFR_X1 \addr_output_reg[18]  (.D(n_0_70), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_0), .QN());
   DFFR_X1 \addr_output_reg[17]  (.D(n_0_69), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_1), .QN());
   DFFR_X1 \addr_output_reg[16]  (.D(n_0_68), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_2), .QN());
   DFFR_X1 \addr_output_reg[15]  (.D(n_0_67), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_36), .QN());
   DFFR_X1 \addr_output_reg[14]  (.D(n_0_66), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_37), .QN());
   DFFR_X1 \addr_output_reg[13]  (.D(n_0_65), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_38), .QN());
   DFFR_X1 \addr_output_reg[12]  (.D(n_0_64), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_39), .QN());
   DFFS_X1 \addr_output_reg[11]  (.D(n_0_63), .SN(n_0_295), .CK(n_0_269), 
      .Q(n_0_40), .QN());
   DFFR_X1 \addr_output_reg[10]  (.D(n_0_62), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_41), .QN());
   DFFR_X1 \addr_output_reg[9]  (.D(n_0_61), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_42), .QN());
   DFFS_X1 \addr_output_reg[8]  (.D(n_0_60), .SN(n_0_295), .CK(n_0_269), 
      .Q(n_0_43), .QN());
   DFFS_X1 \addr_output_reg[7]  (.D(n_0_59), .SN(n_0_295), .CK(n_0_269), 
      .Q(n_0_44), .QN());
   DFFS_X1 \addr_output_reg[6]  (.D(n_0_58), .SN(n_0_295), .CK(n_0_269), 
      .Q(n_0_45), .QN());
   DFFR_X1 \addr_output_reg[5]  (.D(n_0_57), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_46), .QN());
   DFFR_X1 \addr_output_reg[4]  (.D(n_0_56), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_47), .QN());
   DFFR_X1 \addr_output_reg[3]  (.D(n_0_55), .RN(n_0_295), .CK(n_0_269), 
      .Q(n_0_48), .QN());
   DFFS_X1 \addr_output_reg[2]  (.D(n_0_54), .SN(n_0_295), .CK(n_0_269), 
      .Q(n_0_49), .QN());
   DFFS_X1 \addr_output_reg[1]  (.D(n_0_53), .SN(n_0_295), .CK(n_0_269), 
      .Q(n_0_50), .QN());
   DFFS_X1 \addr_output_reg[0]  (.D(n_0_52), .SN(n_0_295), .CK(n_0_269), 
      .Q(n_0_51), .QN());
   datapath__0_144 i_0_18 (.addr_output({n_0_270, n_0_272, n_0_274, n_0_276, 
      n_0_278, n_0_280, n_0_282, n_0_284, n_0_286, n_0_288, n_0_290, n_0_292, 
      n_0_294, n_0_0, n_0_1, n_0_2, n_0_36, n_0_37, n_0_38, n_0_39, n_0_40, 
      n_0_41, n_0_42, n_0_43, n_0_44, n_0_45, n_0_46, n_0_47, n_0_48, n_0_49, 
      n_0_50, n_0_51}), .p_0({n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, 
      n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
      n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, 
      n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52}));
   CLKGATETST_X1 clk_gate_addr_T_reg (.CK(CLK), .E(n_0_118), .SE(1'b0), .GCK(
      n_0_84));
   DFFR_X1 \addr_T_reg[31]  (.D(n_0_35), .RN(n_0_295), .CK(n_0_84), .Q(n_0_85), 
      .QN());
   DFFR_X1 \addr_T_reg[30]  (.D(n_0_34), .RN(n_0_295), .CK(n_0_84), .Q(n_0_86), 
      .QN());
   DFFR_X1 \addr_T_reg[29]  (.D(n_0_33), .RN(n_0_295), .CK(n_0_84), .Q(n_0_87), 
      .QN());
   DFFR_X1 \addr_T_reg[28]  (.D(n_0_32), .RN(n_0_295), .CK(n_0_84), .Q(n_0_88), 
      .QN());
   DFFR_X1 \addr_T_reg[27]  (.D(n_0_31), .RN(n_0_295), .CK(n_0_84), .Q(n_0_89), 
      .QN());
   DFFR_X1 \addr_T_reg[26]  (.D(n_0_30), .RN(n_0_295), .CK(n_0_84), .Q(n_0_90), 
      .QN());
   DFFR_X1 \addr_T_reg[25]  (.D(n_0_29), .RN(n_0_295), .CK(n_0_84), .Q(n_0_91), 
      .QN());
   DFFR_X1 \addr_T_reg[24]  (.D(n_0_28), .RN(n_0_295), .CK(n_0_84), .Q(n_0_92), 
      .QN());
   DFFR_X1 \addr_T_reg[23]  (.D(n_0_27), .RN(n_0_295), .CK(n_0_84), .Q(n_0_93), 
      .QN());
   DFFR_X1 \addr_T_reg[22]  (.D(n_0_26), .RN(n_0_295), .CK(n_0_84), .Q(n_0_94), 
      .QN());
   DFFR_X1 \addr_T_reg[21]  (.D(n_0_25), .RN(n_0_295), .CK(n_0_84), .Q(n_0_95), 
      .QN());
   DFFR_X1 \addr_T_reg[20]  (.D(n_0_24), .RN(n_0_295), .CK(n_0_84), .Q(n_0_96), 
      .QN());
   DFFR_X1 \addr_T_reg[19]  (.D(n_0_23), .RN(n_0_295), .CK(n_0_84), .Q(n_0_97), 
      .QN());
   DFFR_X1 \addr_T_reg[18]  (.D(n_0_22), .RN(n_0_295), .CK(n_0_84), .Q(n_0_98), 
      .QN());
   DFFR_X1 \addr_T_reg[17]  (.D(n_0_21), .RN(n_0_295), .CK(n_0_84), .Q(n_0_99), 
      .QN());
   DFFR_X1 \addr_T_reg[16]  (.D(n_0_20), .RN(n_0_295), .CK(n_0_84), .Q(n_0_100), 
      .QN());
   DFFR_X1 \addr_T_reg[15]  (.D(n_0_19), .RN(n_0_295), .CK(n_0_84), .Q(n_0_101), 
      .QN());
   DFFR_X1 \addr_T_reg[14]  (.D(n_0_18), .RN(n_0_295), .CK(n_0_84), .Q(n_0_102), 
      .QN());
   DFFR_X1 \addr_T_reg[13]  (.D(n_0_17), .RN(n_0_295), .CK(n_0_84), .Q(n_0_103), 
      .QN());
   DFFS_X1 \addr_T_reg[12]  (.D(n_0_16), .SN(n_0_295), .CK(n_0_84), .Q(n_0_104), 
      .QN());
   DFFR_X1 \addr_T_reg[11]  (.D(n_0_15), .RN(n_0_295), .CK(n_0_84), .Q(n_0_105), 
      .QN());
   DFFR_X1 \addr_T_reg[10]  (.D(n_0_14), .RN(n_0_295), .CK(n_0_84), .Q(n_0_106), 
      .QN());
   DFFS_X1 \addr_T_reg[9]  (.D(n_0_13), .SN(n_0_295), .CK(n_0_84), .Q(n_0_107), 
      .QN());
   DFFS_X1 \addr_T_reg[8]  (.D(n_0_12), .SN(n_0_295), .CK(n_0_84), .Q(n_0_108), 
      .QN());
   DFFS_X1 \addr_T_reg[7]  (.D(n_0_11), .SN(n_0_295), .CK(n_0_84), .Q(n_0_109), 
      .QN());
   DFFR_X1 \addr_T_reg[6]  (.D(n_0_10), .RN(n_0_295), .CK(n_0_84), .Q(n_0_110), 
      .QN());
   DFFR_X1 \addr_T_reg[5]  (.D(n_0_9), .RN(n_0_295), .CK(n_0_84), .Q(n_0_111), 
      .QN());
   DFFR_X1 \addr_T_reg[4]  (.D(n_0_8), .RN(n_0_295), .CK(n_0_84), .Q(n_0_112), 
      .QN());
   DFFS_X1 \addr_T_reg[3]  (.D(n_0_7), .SN(n_0_295), .CK(n_0_84), .Q(n_0_113), 
      .QN());
   DFFR_X1 \addr_T_reg[2]  (.D(n_0_6), .RN(n_0_295), .CK(n_0_84), .Q(n_0_114), 
      .QN());
   DFFS_X1 \addr_T_reg[1]  (.D(n_0_5), .SN(n_0_295), .CK(n_0_84), .Q(n_0_115), 
      .QN());
   DFFS_X1 \addr_T_reg[0]  (.D(n_0_4), .SN(n_0_295), .CK(n_0_84), .Q(n_0_116), 
      .QN());
   DFFR_X1 \state_reg[0]__0  (.D(n_0_117), .RN(n_0_295), .CK(n_0_201), .Q(
      state[0]), .QN());
   AND2_X1 i_0_0_0 (.A1(n_0_0_104), .A2(n_0_0_37), .ZN(n_0_119));
   INV_X1 i_0_0_1 (.A(n_0_0_0), .ZN(n_0_232));
   AOI222_X1 i_0_0_2 (.A1(memory_data[0]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[32]), .C1(CPU_Bus[0]), .C2(n_0_0_35), .ZN(n_0_0_0));
   INV_X1 i_0_0_3 (.A(n_0_0_1), .ZN(n_0_231));
   AOI222_X1 i_0_0_4 (.A1(memory_data[1]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[33]), .C1(CPU_Bus[1]), .C2(n_0_0_35), .ZN(n_0_0_1));
   INV_X1 i_0_0_5 (.A(n_0_0_2), .ZN(n_0_230));
   AOI222_X1 i_0_0_6 (.A1(memory_data[2]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[34]), .C1(CPU_Bus[2]), .C2(n_0_0_35), .ZN(n_0_0_2));
   INV_X1 i_0_0_7 (.A(n_0_0_3), .ZN(n_0_229));
   AOI222_X1 i_0_0_8 (.A1(memory_data[3]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[35]), .C1(CPU_Bus[3]), .C2(n_0_0_35), .ZN(n_0_0_3));
   INV_X1 i_0_0_9 (.A(n_0_0_4), .ZN(n_0_228));
   AOI222_X1 i_0_0_10 (.A1(memory_data[4]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[36]), .C1(CPU_Bus[4]), .C2(n_0_0_35), .ZN(n_0_0_4));
   INV_X1 i_0_0_11 (.A(n_0_0_5), .ZN(n_0_227));
   AOI222_X1 i_0_0_12 (.A1(memory_data[5]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[37]), .C1(CPU_Bus[5]), .C2(n_0_0_35), .ZN(n_0_0_5));
   INV_X1 i_0_0_13 (.A(n_0_0_6), .ZN(n_0_226));
   AOI222_X1 i_0_0_14 (.A1(memory_data[6]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[38]), .C1(CPU_Bus[6]), .C2(n_0_0_35), .ZN(n_0_0_6));
   INV_X1 i_0_0_15 (.A(n_0_0_7), .ZN(n_0_225));
   AOI222_X1 i_0_0_16 (.A1(memory_data[7]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[39]), .C1(CPU_Bus[7]), .C2(n_0_0_35), .ZN(n_0_0_7));
   INV_X1 i_0_0_17 (.A(n_0_0_8), .ZN(n_0_224));
   AOI222_X1 i_0_0_18 (.A1(memory_data[8]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[40]), .C1(CPU_Bus[8]), .C2(n_0_0_35), .ZN(n_0_0_8));
   INV_X1 i_0_0_19 (.A(n_0_0_9), .ZN(n_0_223));
   AOI222_X1 i_0_0_20 (.A1(memory_data[9]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[41]), .C1(CPU_Bus[9]), .C2(n_0_0_35), .ZN(n_0_0_9));
   INV_X1 i_0_0_21 (.A(n_0_0_10), .ZN(n_0_222));
   AOI222_X1 i_0_0_22 (.A1(memory_data[10]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[42]), .C1(CPU_Bus[10]), .C2(n_0_0_35), .ZN(n_0_0_10));
   INV_X1 i_0_0_23 (.A(n_0_0_11), .ZN(n_0_221));
   AOI222_X1 i_0_0_24 (.A1(memory_data[11]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[43]), .C1(CPU_Bus[11]), .C2(n_0_0_35), .ZN(n_0_0_11));
   INV_X1 i_0_0_25 (.A(n_0_0_12), .ZN(n_0_220));
   AOI222_X1 i_0_0_26 (.A1(memory_data[12]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[44]), .C1(CPU_Bus[12]), .C2(n_0_0_35), .ZN(n_0_0_12));
   INV_X1 i_0_0_27 (.A(n_0_0_13), .ZN(n_0_219));
   AOI222_X1 i_0_0_28 (.A1(memory_data[13]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[45]), .C1(CPU_Bus[13]), .C2(n_0_0_35), .ZN(n_0_0_13));
   INV_X1 i_0_0_29 (.A(n_0_0_14), .ZN(n_0_218));
   AOI222_X1 i_0_0_30 (.A1(memory_data[14]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[46]), .C1(CPU_Bus[14]), .C2(n_0_0_35), .ZN(n_0_0_14));
   INV_X1 i_0_0_31 (.A(n_0_0_15), .ZN(n_0_217));
   AOI222_X1 i_0_0_32 (.A1(memory_data[15]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[47]), .C1(CPU_Bus[15]), .C2(n_0_0_35), .ZN(n_0_0_15));
   INV_X1 i_0_0_33 (.A(n_0_0_16), .ZN(n_0_216));
   AOI222_X1 i_0_0_34 (.A1(memory_data[16]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[48]), .C1(CPU_Bus[16]), .C2(n_0_0_35), .ZN(n_0_0_16));
   INV_X1 i_0_0_35 (.A(n_0_0_17), .ZN(n_0_215));
   AOI222_X1 i_0_0_36 (.A1(memory_data[17]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[49]), .C1(CPU_Bus[17]), .C2(n_0_0_35), .ZN(n_0_0_17));
   INV_X1 i_0_0_37 (.A(n_0_0_18), .ZN(n_0_214));
   AOI222_X1 i_0_0_38 (.A1(memory_data[18]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[50]), .C1(CPU_Bus[18]), .C2(n_0_0_35), .ZN(n_0_0_18));
   INV_X1 i_0_0_39 (.A(n_0_0_19), .ZN(n_0_213));
   AOI222_X1 i_0_0_40 (.A1(memory_data[19]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[51]), .C1(CPU_Bus[19]), .C2(n_0_0_35), .ZN(n_0_0_19));
   INV_X1 i_0_0_41 (.A(n_0_0_20), .ZN(n_0_212));
   AOI222_X1 i_0_0_42 (.A1(memory_data[20]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[52]), .C1(CPU_Bus[20]), .C2(n_0_0_35), .ZN(n_0_0_20));
   INV_X1 i_0_0_43 (.A(n_0_0_21), .ZN(n_0_211));
   AOI222_X1 i_0_0_44 (.A1(memory_data[21]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[53]), .C1(CPU_Bus[21]), .C2(n_0_0_35), .ZN(n_0_0_21));
   INV_X1 i_0_0_45 (.A(n_0_0_22), .ZN(n_0_210));
   AOI222_X1 i_0_0_46 (.A1(memory_data[22]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[54]), .C1(CPU_Bus[22]), .C2(n_0_0_35), .ZN(n_0_0_22));
   INV_X1 i_0_0_47 (.A(n_0_0_23), .ZN(n_0_209));
   AOI222_X1 i_0_0_48 (.A1(memory_data[23]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[55]), .C1(CPU_Bus[23]), .C2(n_0_0_35), .ZN(n_0_0_23));
   INV_X1 i_0_0_49 (.A(n_0_0_24), .ZN(n_0_208));
   AOI222_X1 i_0_0_50 (.A1(memory_data[24]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[56]), .C1(CPU_Bus[24]), .C2(n_0_0_35), .ZN(n_0_0_24));
   INV_X1 i_0_0_51 (.A(n_0_0_25), .ZN(n_0_207));
   AOI222_X1 i_0_0_52 (.A1(memory_data[25]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[57]), .C1(CPU_Bus[25]), .C2(n_0_0_35), .ZN(n_0_0_25));
   INV_X1 i_0_0_53 (.A(n_0_0_26), .ZN(n_0_206));
   AOI222_X1 i_0_0_54 (.A1(memory_data[26]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[58]), .C1(CPU_Bus[26]), .C2(n_0_0_35), .ZN(n_0_0_26));
   INV_X1 i_0_0_55 (.A(n_0_0_27), .ZN(n_0_205));
   AOI222_X1 i_0_0_56 (.A1(memory_data[27]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[59]), .C1(CPU_Bus[27]), .C2(n_0_0_35), .ZN(n_0_0_27));
   INV_X1 i_0_0_57 (.A(n_0_0_28), .ZN(n_0_204));
   AOI222_X1 i_0_0_58 (.A1(memory_data[28]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[60]), .C1(CPU_Bus[28]), .C2(n_0_0_35), .ZN(n_0_0_28));
   INV_X1 i_0_0_59 (.A(n_0_0_29), .ZN(n_0_203));
   AOI222_X1 i_0_0_60 (.A1(memory_data[29]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[61]), .C1(CPU_Bus[29]), .C2(n_0_0_35), .ZN(n_0_0_29));
   INV_X1 i_0_0_61 (.A(n_0_0_30), .ZN(n_0_202));
   AOI222_X1 i_0_0_62 (.A1(memory_data[30]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[62]), .C1(CPU_Bus[30]), .C2(n_0_0_35), .ZN(n_0_0_30));
   INV_X1 i_0_0_63 (.A(n_0_0_31), .ZN(n_0_200));
   AOI222_X1 i_0_0_64 (.A1(memory_data[31]), .A2(n_0_0_33), .B1(n_0_0_32), 
      .B2(memory_data[63]), .C1(CPU_Bus[31]), .C2(n_0_0_35), .ZN(n_0_0_31));
   NOR3_X1 i_0_0_65 (.A1(n_0_0_35), .A2(state_reg[0]), .A3(state_reg[1]), 
      .ZN(n_0_0_32));
   AOI21_X1 i_0_0_66 (.A(n_0_0_35), .B1(n_0_117), .B2(n_0_0_34), .ZN(n_0_0_33));
   OR2_X1 i_0_0_67 (.A1(n_0_0_158), .A2(state_reg[0]), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_68 (.A1(n_0_0_158), .A2(state_reg[0]), .ZN(n_0_117));
   NAND2_X1 i_0_0_69 (.A1(n_0_0_159), .A2(enable_output_IO), .ZN(n_0_0_35));
   AND2_X1 i_0_0_70 (.A1(n_0_0_36), .A2(memory_address[0]), .ZN(n_0_198));
   AND2_X1 i_0_0_71 (.A1(n_0_0_36), .A2(memory_address[1]), .ZN(n_0_197));
   AND2_X1 i_0_0_72 (.A1(n_0_0_36), .A2(memory_address[2]), .ZN(n_0_196));
   AND2_X1 i_0_0_73 (.A1(n_0_0_36), .A2(memory_address[3]), .ZN(n_0_195));
   AND2_X1 i_0_0_74 (.A1(n_0_0_36), .A2(memory_address[4]), .ZN(n_0_194));
   AND2_X1 i_0_0_75 (.A1(n_0_0_36), .A2(memory_address[5]), .ZN(n_0_193));
   AND2_X1 i_0_0_76 (.A1(n_0_0_36), .A2(memory_address[6]), .ZN(n_0_192));
   AND2_X1 i_0_0_77 (.A1(n_0_0_36), .A2(memory_address[7]), .ZN(n_0_191));
   AND2_X1 i_0_0_78 (.A1(n_0_0_36), .A2(memory_address[8]), .ZN(n_0_190));
   AND2_X1 i_0_0_79 (.A1(n_0_0_36), .A2(memory_address[9]), .ZN(n_0_189));
   AND2_X1 i_0_0_80 (.A1(n_0_0_36), .A2(memory_address[10]), .ZN(n_0_188));
   AND2_X1 i_0_0_81 (.A1(n_0_0_36), .A2(memory_address[11]), .ZN(n_0_187));
   AND2_X1 i_0_0_82 (.A1(n_0_0_36), .A2(memory_address[12]), .ZN(n_0_186));
   AND2_X1 i_0_0_83 (.A1(n_0_0_36), .A2(memory_address[13]), .ZN(n_0_185));
   AND2_X1 i_0_0_84 (.A1(n_0_0_36), .A2(memory_address[14]), .ZN(n_0_184));
   AND2_X1 i_0_0_85 (.A1(n_0_0_36), .A2(memory_address[15]), .ZN(n_0_183));
   AND2_X1 i_0_0_86 (.A1(n_0_0_36), .A2(memory_address[16]), .ZN(n_0_182));
   AND2_X1 i_0_0_87 (.A1(n_0_0_36), .A2(memory_address[17]), .ZN(n_0_181));
   AND2_X1 i_0_0_88 (.A1(n_0_0_36), .A2(memory_address[18]), .ZN(n_0_180));
   AND2_X1 i_0_0_89 (.A1(n_0_0_36), .A2(memory_address[19]), .ZN(n_0_179));
   AND2_X1 i_0_0_90 (.A1(n_0_0_36), .A2(memory_address[20]), .ZN(n_0_178));
   AND2_X1 i_0_0_91 (.A1(n_0_0_36), .A2(memory_address[21]), .ZN(n_0_177));
   AND2_X1 i_0_0_92 (.A1(n_0_0_36), .A2(memory_address[22]), .ZN(n_0_176));
   AND2_X1 i_0_0_93 (.A1(n_0_0_36), .A2(memory_address[23]), .ZN(n_0_175));
   AND2_X1 i_0_0_94 (.A1(n_0_0_36), .A2(memory_address[24]), .ZN(n_0_174));
   AND2_X1 i_0_0_95 (.A1(n_0_0_36), .A2(memory_address[25]), .ZN(n_0_173));
   AND2_X1 i_0_0_96 (.A1(n_0_0_36), .A2(memory_address[26]), .ZN(n_0_172));
   AND2_X1 i_0_0_97 (.A1(n_0_0_36), .A2(memory_address[27]), .ZN(n_0_171));
   AND2_X1 i_0_0_98 (.A1(n_0_0_36), .A2(memory_address[28]), .ZN(n_0_170));
   AND2_X1 i_0_0_99 (.A1(n_0_0_36), .A2(memory_address[29]), .ZN(n_0_169));
   AND2_X1 i_0_0_100 (.A1(n_0_0_36), .A2(memory_address[30]), .ZN(n_0_168));
   AND2_X1 i_0_0_101 (.A1(n_0_0_36), .A2(memory_address[31]), .ZN(n_0_167));
   NAND3_X1 i_0_0_102 (.A1(enable_output_IO), .A2(state_reg[1]), .A3(
      state_reg[0]), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_103 (.A1(n_0_116), .A2(RST), .ZN(n_0_135));
   NAND2_X1 i_0_0_104 (.A1(n_0_115), .A2(RST), .ZN(n_0_136));
   NAND2_X1 i_0_0_105 (.A1(n_0_114), .A2(RST), .ZN(n_0_137));
   NAND2_X1 i_0_0_106 (.A1(n_0_113), .A2(RST), .ZN(n_0_138));
   NAND2_X1 i_0_0_107 (.A1(n_0_112), .A2(RST), .ZN(n_0_139));
   NAND2_X1 i_0_0_108 (.A1(n_0_111), .A2(RST), .ZN(n_0_140));
   NAND2_X1 i_0_0_109 (.A1(n_0_110), .A2(RST), .ZN(n_0_141));
   NAND2_X1 i_0_0_110 (.A1(n_0_109), .A2(RST), .ZN(n_0_142));
   NAND2_X1 i_0_0_111 (.A1(n_0_108), .A2(RST), .ZN(n_0_143));
   NAND2_X1 i_0_0_112 (.A1(n_0_107), .A2(RST), .ZN(n_0_144));
   NAND2_X1 i_0_0_113 (.A1(n_0_106), .A2(RST), .ZN(n_0_145));
   NAND2_X1 i_0_0_114 (.A1(n_0_105), .A2(RST), .ZN(n_0_146));
   NAND2_X1 i_0_0_115 (.A1(n_0_104), .A2(RST), .ZN(n_0_147));
   NAND2_X1 i_0_0_116 (.A1(n_0_103), .A2(RST), .ZN(n_0_148));
   NAND2_X1 i_0_0_117 (.A1(n_0_102), .A2(RST), .ZN(n_0_149));
   NAND2_X1 i_0_0_118 (.A1(n_0_101), .A2(RST), .ZN(n_0_150));
   NAND2_X1 i_0_0_119 (.A1(n_0_100), .A2(RST), .ZN(n_0_151));
   NAND2_X1 i_0_0_120 (.A1(n_0_99), .A2(RST), .ZN(n_0_152));
   NAND2_X1 i_0_0_121 (.A1(n_0_98), .A2(RST), .ZN(n_0_153));
   NAND2_X1 i_0_0_122 (.A1(n_0_97), .A2(RST), .ZN(n_0_154));
   NAND2_X1 i_0_0_123 (.A1(n_0_96), .A2(RST), .ZN(n_0_155));
   NAND2_X1 i_0_0_124 (.A1(n_0_95), .A2(RST), .ZN(n_0_156));
   NAND2_X1 i_0_0_125 (.A1(n_0_94), .A2(RST), .ZN(n_0_157));
   NAND2_X1 i_0_0_126 (.A1(n_0_93), .A2(RST), .ZN(n_0_158));
   NAND2_X1 i_0_0_127 (.A1(n_0_92), .A2(RST), .ZN(n_0_159));
   NAND2_X1 i_0_0_128 (.A1(n_0_91), .A2(RST), .ZN(n_0_160));
   NAND2_X1 i_0_0_129 (.A1(n_0_90), .A2(RST), .ZN(n_0_161));
   NAND2_X1 i_0_0_130 (.A1(n_0_89), .A2(RST), .ZN(n_0_162));
   NAND2_X1 i_0_0_131 (.A1(n_0_88), .A2(RST), .ZN(n_0_163));
   NAND2_X1 i_0_0_132 (.A1(n_0_87), .A2(RST), .ZN(n_0_164));
   NAND2_X1 i_0_0_133 (.A1(n_0_86), .A2(RST), .ZN(n_0_165));
   NAND2_X1 i_0_0_134 (.A1(n_0_85), .A2(RST), .ZN(n_0_166));
   NAND2_X1 i_0_0_135 (.A1(n_0_0_191), .A2(RST), .ZN(n_0_120));
   NAND2_X1 i_0_0_136 (.A1(n_0_0_192), .A2(RST), .ZN(n_0_121));
   NAND2_X1 i_0_0_137 (.A1(n_0_0_193), .A2(RST), .ZN(n_0_122));
   NAND2_X1 i_0_0_138 (.A1(n_0_0_194), .A2(RST), .ZN(n_0_123));
   NAND2_X1 i_0_0_139 (.A1(n_0_0_195), .A2(RST), .ZN(n_0_124));
   NAND2_X1 i_0_0_140 (.A1(n_0_0_196), .A2(RST), .ZN(n_0_125));
   NAND2_X1 i_0_0_141 (.A1(n_0_0_197), .A2(RST), .ZN(n_0_126));
   NAND2_X1 i_0_0_142 (.A1(n_0_0_198), .A2(RST), .ZN(n_0_127));
   NAND2_X1 i_0_0_143 (.A1(n_0_0_199), .A2(RST), .ZN(n_0_128));
   NAND2_X1 i_0_0_144 (.A1(n_0_0_200), .A2(RST), .ZN(n_0_129));
   NAND2_X1 i_0_0_145 (.A1(n_0_0_201), .A2(RST), .ZN(n_0_130));
   NAND2_X1 i_0_0_146 (.A1(n_0_0_202), .A2(RST), .ZN(n_0_131));
   NAND2_X1 i_0_0_147 (.A1(n_0_0_203), .A2(RST), .ZN(n_0_132));
   NAND2_X1 i_0_0_148 (.A1(n_0_0_204), .A2(RST), .ZN(n_0_133));
   NAND2_X1 i_0_0_149 (.A1(n_0_0_205), .A2(RST), .ZN(n_0_134));
   NAND2_X1 i_0_0_150 (.A1(n_0_0_206), .A2(RST), .ZN(n_0_199));
   NAND2_X1 i_0_0_151 (.A1(n_0_0_207), .A2(RST), .ZN(n_0_233));
   NAND2_X1 i_0_0_152 (.A1(n_0_0_208), .A2(RST), .ZN(n_0_234));
   NAND2_X1 i_0_0_153 (.A1(n_0_0_209), .A2(RST), .ZN(n_0_235));
   NAND2_X1 i_0_0_154 (.A1(n_0_0_210), .A2(RST), .ZN(n_0_236));
   NAND2_X1 i_0_0_155 (.A1(n_0_0_211), .A2(RST), .ZN(n_0_237));
   NAND2_X1 i_0_0_156 (.A1(n_0_0_212), .A2(RST), .ZN(n_0_238));
   NAND2_X1 i_0_0_157 (.A1(n_0_0_213), .A2(RST), .ZN(n_0_239));
   NAND2_X1 i_0_0_158 (.A1(n_0_0_214), .A2(RST), .ZN(n_0_240));
   NAND2_X1 i_0_0_159 (.A1(n_0_0_215), .A2(RST), .ZN(n_0_241));
   NAND2_X1 i_0_0_160 (.A1(n_0_0_216), .A2(RST), .ZN(n_0_242));
   NAND2_X1 i_0_0_161 (.A1(n_0_0_217), .A2(RST), .ZN(n_0_243));
   NAND2_X1 i_0_0_162 (.A1(n_0_0_218), .A2(RST), .ZN(n_0_244));
   NAND2_X1 i_0_0_163 (.A1(n_0_0_219), .A2(RST), .ZN(n_0_245));
   NAND2_X1 i_0_0_164 (.A1(n_0_0_220), .A2(RST), .ZN(n_0_246));
   NAND2_X1 i_0_0_165 (.A1(n_0_0_221), .A2(RST), .ZN(n_0_247));
   OR2_X1 i_0_0_166 (.A1(n_0_0_159), .A2(n_0_85), .ZN(n_0_248));
   OR2_X1 i_0_0_167 (.A1(n_0_118), .A2(n_0_0_37), .ZN(eq));
   NOR3_X1 i_0_0_168 (.A1(done_output_data), .A2(state[0]), .A3(n_0_0_38), 
      .ZN(n_0_0_37));
   AOI21_X1 i_0_0_169 (.A(n_0_0_39), .B1(n_0_270), .B2(n_0_0_190), .ZN(n_0_0_38));
   NOR2_X1 i_0_0_170 (.A1(n_0_0_41), .A2(n_0_0_40), .ZN(n_0_0_39));
   OAI22_X1 i_0_0_171 (.A1(n_0_0_190), .A2(n_0_270), .B1(n_0_0_174), .B2(
      end_Output_address[30]), .ZN(n_0_0_40));
   AOI21_X1 i_0_0_172 (.A(n_0_0_42), .B1(n_0_0_174), .B2(end_Output_address[30]), 
      .ZN(n_0_0_41));
   AOI21_X1 i_0_0_173 (.A(n_0_0_86), .B1(n_0_0_44), .B2(n_0_0_43), .ZN(n_0_0_42));
   AOI22_X1 i_0_0_174 (.A1(end_Output_address[29]), .A2(n_0_0_173), .B1(
      n_0_0_172), .B2(end_Output_address[28]), .ZN(n_0_0_43));
   OAI221_X1 i_0_0_175 (.A(n_0_0_45), .B1(end_Output_address[28]), .B2(n_0_0_172), 
      .C1(n_0_0_47), .C2(n_0_0_46), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_176 (.A1(n_0_0_189), .A2(n_0_278), .ZN(n_0_0_45));
   OAI22_X1 i_0_0_177 (.A1(n_0_0_189), .A2(n_0_278), .B1(n_0_0_188), .B2(n_0_280), 
      .ZN(n_0_0_46));
   AOI221_X1 i_0_0_178 (.A(n_0_0_48), .B1(n_0_0_188), .B2(n_0_280), .C1(n_0_0_50), 
      .C2(n_0_0_49), .ZN(n_0_0_47));
   NOR2_X1 i_0_0_179 (.A1(n_0_0_171), .A2(end_Output_address[25]), .ZN(n_0_0_48));
   AOI22_X1 i_0_0_180 (.A1(end_Output_address[25]), .A2(n_0_0_171), .B1(
      n_0_0_170), .B2(end_Output_address[24]), .ZN(n_0_0_49));
   OAI221_X1 i_0_0_181 (.A(n_0_0_51), .B1(end_Output_address[24]), .B2(n_0_0_170), 
      .C1(n_0_0_53), .C2(n_0_0_52), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_182 (.A1(n_0_0_187), .A2(n_0_286), .ZN(n_0_0_51));
   OAI22_X1 i_0_0_183 (.A1(n_0_0_187), .A2(n_0_286), .B1(n_0_0_186), .B2(n_0_288), 
      .ZN(n_0_0_52));
   AOI221_X1 i_0_0_184 (.A(n_0_0_54), .B1(n_0_0_186), .B2(n_0_288), .C1(n_0_0_56), 
      .C2(n_0_0_55), .ZN(n_0_0_53));
   NOR2_X1 i_0_0_185 (.A1(n_0_0_169), .A2(end_Output_address[21]), .ZN(n_0_0_54));
   AOI22_X1 i_0_0_186 (.A1(end_Output_address[21]), .A2(n_0_0_169), .B1(
      n_0_0_168), .B2(end_Output_address[20]), .ZN(n_0_0_55));
   OAI221_X1 i_0_0_187 (.A(n_0_0_57), .B1(end_Output_address[20]), .B2(n_0_0_168), 
      .C1(n_0_0_59), .C2(n_0_0_58), .ZN(n_0_0_56));
   NAND2_X1 i_0_0_188 (.A1(n_0_0_185), .A2(n_0_294), .ZN(n_0_0_57));
   OAI22_X1 i_0_0_189 (.A1(n_0_0_185), .A2(n_0_294), .B1(n_0_0_184), .B2(n_0_0), 
      .ZN(n_0_0_58));
   AOI221_X1 i_0_0_190 (.A(n_0_0_60), .B1(n_0_0_184), .B2(n_0_0), .C1(n_0_0_62), 
      .C2(n_0_0_61), .ZN(n_0_0_59));
   NOR2_X1 i_0_0_191 (.A1(n_0_0_167), .A2(end_Output_address[17]), .ZN(n_0_0_60));
   AOI22_X1 i_0_0_192 (.A1(end_Output_address[17]), .A2(n_0_0_167), .B1(
      n_0_0_166), .B2(end_Output_address[16]), .ZN(n_0_0_61));
   OAI221_X1 i_0_0_193 (.A(n_0_0_63), .B1(end_Output_address[16]), .B2(n_0_0_166), 
      .C1(n_0_0_65), .C2(n_0_0_64), .ZN(n_0_0_62));
   NAND2_X1 i_0_0_194 (.A1(n_0_0_183), .A2(n_0_36), .ZN(n_0_0_63));
   OAI22_X1 i_0_0_195 (.A1(n_0_0_183), .A2(n_0_36), .B1(n_0_0_182), .B2(n_0_37), 
      .ZN(n_0_0_64));
   AOI221_X1 i_0_0_196 (.A(n_0_0_66), .B1(n_0_0_182), .B2(n_0_37), .C1(n_0_0_68), 
      .C2(n_0_0_67), .ZN(n_0_0_65));
   NOR2_X1 i_0_0_197 (.A1(n_0_0_165), .A2(end_Output_address[13]), .ZN(n_0_0_66));
   AOI22_X1 i_0_0_198 (.A1(end_Output_address[13]), .A2(n_0_0_165), .B1(
      n_0_0_164), .B2(end_Output_address[12]), .ZN(n_0_0_67));
   OAI221_X1 i_0_0_199 (.A(n_0_0_69), .B1(end_Output_address[12]), .B2(n_0_0_164), 
      .C1(n_0_0_71), .C2(n_0_0_70), .ZN(n_0_0_68));
   NAND2_X1 i_0_0_200 (.A1(n_0_0_181), .A2(n_0_40), .ZN(n_0_0_69));
   OAI22_X1 i_0_0_201 (.A1(n_0_0_181), .A2(n_0_40), .B1(n_0_0_180), .B2(n_0_41), 
      .ZN(n_0_0_70));
   AOI221_X1 i_0_0_202 (.A(n_0_0_72), .B1(n_0_0_180), .B2(n_0_41), .C1(n_0_0_74), 
      .C2(n_0_0_73), .ZN(n_0_0_71));
   NOR2_X1 i_0_0_203 (.A1(n_0_0_163), .A2(end_Output_address[9]), .ZN(n_0_0_72));
   AOI22_X1 i_0_0_204 (.A1(end_Output_address[9]), .A2(n_0_0_163), .B1(n_0_0_162), 
      .B2(end_Output_address[8]), .ZN(n_0_0_73));
   OAI221_X1 i_0_0_205 (.A(n_0_0_75), .B1(end_Output_address[8]), .B2(n_0_0_162), 
      .C1(n_0_0_77), .C2(n_0_0_76), .ZN(n_0_0_74));
   NAND2_X1 i_0_0_206 (.A1(n_0_0_179), .A2(n_0_44), .ZN(n_0_0_75));
   OAI22_X1 i_0_0_207 (.A1(n_0_0_179), .A2(n_0_44), .B1(n_0_0_178), .B2(n_0_45), 
      .ZN(n_0_0_76));
   AOI221_X1 i_0_0_208 (.A(n_0_0_78), .B1(n_0_0_178), .B2(n_0_45), .C1(n_0_0_80), 
      .C2(n_0_0_79), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_209 (.A1(n_0_0_161), .A2(end_Output_address[5]), .ZN(n_0_0_78));
   AOI22_X1 i_0_0_210 (.A1(end_Output_address[5]), .A2(n_0_0_161), .B1(n_0_0_160), 
      .B2(end_Output_address[4]), .ZN(n_0_0_79));
   OAI221_X1 i_0_0_211 (.A(n_0_0_81), .B1(end_Output_address[4]), .B2(n_0_0_160), 
      .C1(n_0_0_83), .C2(n_0_0_82), .ZN(n_0_0_80));
   NAND2_X1 i_0_0_212 (.A1(n_0_0_177), .A2(n_0_48), .ZN(n_0_0_81));
   OAI22_X1 i_0_0_213 (.A1(n_0_0_177), .A2(n_0_48), .B1(n_0_0_176), .B2(n_0_49), 
      .ZN(n_0_0_82));
   AOI221_X1 i_0_0_214 (.A(n_0_0_84), .B1(n_0_50), .B2(n_0_0_175), .C1(n_0_0_176), 
      .C2(n_0_49), .ZN(n_0_0_83));
   NOR2_X1 i_0_0_215 (.A1(n_0_0_85), .A2(end_Output_address[0]), .ZN(n_0_0_84));
   OAI21_X1 i_0_0_216 (.A(n_0_51), .B1(n_0_0_175), .B2(n_0_50), .ZN(n_0_0_85));
   NOR2_X1 i_0_0_217 (.A1(n_0_0_173), .A2(end_Output_address[29]), .ZN(n_0_0_86));
   OAI21_X1 i_0_0_218 (.A(n_0_0_87), .B1(n_0_0_103), .B2(n_0_116), .ZN(n_0_249));
   NAND2_X1 i_0_0_219 (.A1(n_0_0_103), .A2(n_0_51), .ZN(n_0_0_87));
   MUX2_X1 i_0_0_220 (.A(n_0_5), .B(n_0_50), .S(n_0_0_103), .Z(n_0_250));
   MUX2_X1 i_0_0_221 (.A(n_0_6), .B(n_0_49), .S(n_0_0_103), .Z(n_0_251));
   MUX2_X1 i_0_0_222 (.A(n_0_7), .B(n_0_48), .S(n_0_0_103), .Z(n_0_252));
   OAI21_X1 i_0_0_223 (.A(n_0_0_88), .B1(n_0_118), .B2(n_0_0_160), .ZN(n_0_253));
   NAND2_X1 i_0_0_224 (.A1(n_0_8), .A2(n_0_118), .ZN(n_0_0_88));
   OAI21_X1 i_0_0_225 (.A(n_0_0_89), .B1(n_0_118), .B2(n_0_0_161), .ZN(n_0_254));
   NAND2_X1 i_0_0_226 (.A1(n_0_9), .A2(n_0_118), .ZN(n_0_0_89));
   MUX2_X1 i_0_0_227 (.A(n_0_10), .B(n_0_45), .S(n_0_0_103), .Z(n_0_255));
   MUX2_X1 i_0_0_228 (.A(n_0_11), .B(n_0_44), .S(n_0_0_103), .Z(n_0_256));
   OAI21_X1 i_0_0_229 (.A(n_0_0_90), .B1(n_0_118), .B2(n_0_0_162), .ZN(n_0_257));
   NAND2_X1 i_0_0_230 (.A1(n_0_12), .A2(n_0_118), .ZN(n_0_0_90));
   OAI21_X1 i_0_0_231 (.A(n_0_0_91), .B1(n_0_118), .B2(n_0_0_163), .ZN(n_0_258));
   NAND2_X1 i_0_0_232 (.A1(n_0_13), .A2(n_0_118), .ZN(n_0_0_91));
   MUX2_X1 i_0_0_233 (.A(n_0_14), .B(n_0_41), .S(n_0_0_103), .Z(n_0_259));
   MUX2_X1 i_0_0_234 (.A(n_0_15), .B(n_0_40), .S(n_0_0_103), .Z(n_0_260));
   OAI21_X1 i_0_0_235 (.A(n_0_0_92), .B1(n_0_118), .B2(n_0_0_164), .ZN(n_0_261));
   NAND2_X1 i_0_0_236 (.A1(n_0_16), .A2(n_0_118), .ZN(n_0_0_92));
   OAI21_X1 i_0_0_237 (.A(n_0_0_93), .B1(n_0_118), .B2(n_0_0_165), .ZN(n_0_262));
   NAND2_X1 i_0_0_238 (.A1(n_0_17), .A2(n_0_118), .ZN(n_0_0_93));
   MUX2_X1 i_0_0_239 (.A(n_0_18), .B(n_0_37), .S(n_0_0_103), .Z(n_0_263));
   MUX2_X1 i_0_0_240 (.A(n_0_19), .B(n_0_36), .S(n_0_0_103), .Z(n_0_264));
   OAI21_X1 i_0_0_241 (.A(n_0_0_94), .B1(n_0_118), .B2(n_0_0_166), .ZN(n_0_265));
   NAND2_X1 i_0_0_242 (.A1(n_0_20), .A2(n_0_118), .ZN(n_0_0_94));
   OAI21_X1 i_0_0_243 (.A(n_0_0_95), .B1(n_0_118), .B2(n_0_0_167), .ZN(n_0_266));
   NAND2_X1 i_0_0_244 (.A1(n_0_21), .A2(n_0_118), .ZN(n_0_0_95));
   MUX2_X1 i_0_0_245 (.A(n_0_22), .B(n_0_0), .S(n_0_0_103), .Z(n_0_267));
   MUX2_X1 i_0_0_246 (.A(n_0_23), .B(n_0_294), .S(n_0_0_103), .Z(n_0_268));
   OAI21_X1 i_0_0_247 (.A(n_0_0_96), .B1(n_0_118), .B2(n_0_0_168), .ZN(n_0_271));
   NAND2_X1 i_0_0_248 (.A1(n_0_24), .A2(n_0_118), .ZN(n_0_0_96));
   OAI21_X1 i_0_0_249 (.A(n_0_0_97), .B1(n_0_118), .B2(n_0_0_169), .ZN(n_0_273));
   NAND2_X1 i_0_0_250 (.A1(n_0_25), .A2(n_0_118), .ZN(n_0_0_97));
   MUX2_X1 i_0_0_251 (.A(n_0_26), .B(n_0_288), .S(n_0_0_103), .Z(n_0_275));
   MUX2_X1 i_0_0_252 (.A(n_0_27), .B(n_0_286), .S(n_0_0_103), .Z(n_0_277));
   OAI21_X1 i_0_0_253 (.A(n_0_0_98), .B1(n_0_118), .B2(n_0_0_170), .ZN(n_0_279));
   NAND2_X1 i_0_0_254 (.A1(n_0_28), .A2(n_0_118), .ZN(n_0_0_98));
   OAI21_X1 i_0_0_255 (.A(n_0_0_99), .B1(n_0_118), .B2(n_0_0_171), .ZN(n_0_281));
   NAND2_X1 i_0_0_256 (.A1(n_0_29), .A2(n_0_118), .ZN(n_0_0_99));
   MUX2_X1 i_0_0_257 (.A(n_0_30), .B(n_0_280), .S(n_0_0_103), .Z(n_0_283));
   MUX2_X1 i_0_0_258 (.A(n_0_31), .B(n_0_278), .S(n_0_0_103), .Z(n_0_285));
   OAI21_X1 i_0_0_259 (.A(n_0_0_100), .B1(n_0_118), .B2(n_0_0_172), .ZN(n_0_287));
   NAND2_X1 i_0_0_260 (.A1(n_0_32), .A2(n_0_118), .ZN(n_0_0_100));
   OAI21_X1 i_0_0_261 (.A(n_0_0_101), .B1(n_0_118), .B2(n_0_0_173), .ZN(n_0_289));
   NAND2_X1 i_0_0_262 (.A1(n_0_33), .A2(n_0_118), .ZN(n_0_0_101));
   OAI21_X1 i_0_0_263 (.A(n_0_0_102), .B1(n_0_118), .B2(n_0_0_174), .ZN(n_0_291));
   NAND2_X1 i_0_0_264 (.A1(n_0_34), .A2(n_0_118), .ZN(n_0_0_102));
   MUX2_X1 i_0_0_265 (.A(n_0_35), .B(n_0_270), .S(n_0_0_103), .Z(n_0_293));
   INV_X1 i_0_0_266 (.A(n_0_0_103), .ZN(n_0_118));
   OR3_X1 i_0_0_267 (.A1(n_0_0_104), .A2(state[0]), .A3(done_output_data), 
      .ZN(n_0_0_103));
   OAI21_X1 i_0_0_268 (.A(n_0_0_105), .B1(n_0_85), .B2(n_0_0_222), .ZN(n_0_0_104));
   NAND2_X1 i_0_0_269 (.A1(n_0_0_107), .A2(n_0_0_106), .ZN(n_0_0_105));
   AOI22_X1 i_0_0_270 (.A1(n_0_0_222), .A2(n_0_85), .B1(n_0_0_221), .B2(
      end_T_address[30]), .ZN(n_0_0_106));
   OAI21_X1 i_0_0_271 (.A(n_0_0_108), .B1(n_0_0_220), .B2(end_T_address[29]), 
      .ZN(n_0_0_107));
   AOI21_X1 i_0_0_272 (.A(n_0_0_109), .B1(n_0_0_111), .B2(n_0_0_110), .ZN(
      n_0_0_108));
   NOR2_X1 i_0_0_273 (.A1(n_0_0_221), .A2(end_T_address[30]), .ZN(n_0_0_109));
   AOI22_X1 i_0_0_274 (.A1(end_T_address[29]), .A2(n_0_0_220), .B1(n_0_0_219), 
      .B2(end_T_address[28]), .ZN(n_0_0_110));
   OAI21_X1 i_0_0_275 (.A(n_0_0_112), .B1(n_0_0_218), .B2(end_T_address[27]), 
      .ZN(n_0_0_111));
   AOI21_X1 i_0_0_276 (.A(n_0_0_113), .B1(n_0_0_115), .B2(n_0_0_114), .ZN(
      n_0_0_112));
   NOR2_X1 i_0_0_277 (.A1(n_0_0_219), .A2(end_T_address[28]), .ZN(n_0_0_113));
   AOI22_X1 i_0_0_278 (.A1(end_T_address[27]), .A2(n_0_0_218), .B1(n_0_0_217), 
      .B2(end_T_address[26]), .ZN(n_0_0_114));
   OAI221_X1 i_0_0_279 (.A(n_0_0_116), .B1(n_0_0_216), .B2(end_T_address[25]), 
      .C1(end_T_address[26]), .C2(n_0_0_217), .ZN(n_0_0_115));
   NAND2_X1 i_0_0_280 (.A1(n_0_0_118), .A2(n_0_0_117), .ZN(n_0_0_116));
   AOI22_X1 i_0_0_281 (.A1(end_T_address[25]), .A2(n_0_0_216), .B1(n_0_0_215), 
      .B2(end_T_address[24]), .ZN(n_0_0_117));
   OAI21_X1 i_0_0_282 (.A(n_0_0_119), .B1(n_0_0_214), .B2(end_T_address[23]), 
      .ZN(n_0_0_118));
   AOI21_X1 i_0_0_283 (.A(n_0_0_120), .B1(n_0_0_122), .B2(n_0_0_121), .ZN(
      n_0_0_119));
   NOR2_X1 i_0_0_284 (.A1(n_0_0_215), .A2(end_T_address[24]), .ZN(n_0_0_120));
   AOI22_X1 i_0_0_285 (.A1(end_T_address[23]), .A2(n_0_0_214), .B1(n_0_0_213), 
      .B2(end_T_address[22]), .ZN(n_0_0_121));
   OAI221_X1 i_0_0_286 (.A(n_0_0_123), .B1(n_0_0_212), .B2(end_T_address[21]), 
      .C1(end_T_address[22]), .C2(n_0_0_213), .ZN(n_0_0_122));
   NAND2_X1 i_0_0_287 (.A1(n_0_0_125), .A2(n_0_0_124), .ZN(n_0_0_123));
   AOI22_X1 i_0_0_288 (.A1(end_T_address[21]), .A2(n_0_0_212), .B1(n_0_0_211), 
      .B2(end_T_address[20]), .ZN(n_0_0_124));
   OAI21_X1 i_0_0_289 (.A(n_0_0_126), .B1(n_0_0_210), .B2(end_T_address[19]), 
      .ZN(n_0_0_125));
   AOI21_X1 i_0_0_290 (.A(n_0_0_127), .B1(n_0_0_129), .B2(n_0_0_128), .ZN(
      n_0_0_126));
   NOR2_X1 i_0_0_291 (.A1(n_0_0_211), .A2(end_T_address[20]), .ZN(n_0_0_127));
   AOI22_X1 i_0_0_292 (.A1(end_T_address[19]), .A2(n_0_0_210), .B1(n_0_0_209), 
      .B2(end_T_address[18]), .ZN(n_0_0_128));
   OAI221_X1 i_0_0_293 (.A(n_0_0_130), .B1(n_0_0_208), .B2(end_T_address[17]), 
      .C1(end_T_address[18]), .C2(n_0_0_209), .ZN(n_0_0_129));
   NAND2_X1 i_0_0_294 (.A1(n_0_0_132), .A2(n_0_0_131), .ZN(n_0_0_130));
   AOI22_X1 i_0_0_295 (.A1(end_T_address[17]), .A2(n_0_0_208), .B1(n_0_0_207), 
      .B2(end_T_address[16]), .ZN(n_0_0_131));
   OAI21_X1 i_0_0_296 (.A(n_0_0_133), .B1(n_0_0_207), .B2(end_T_address[16]), 
      .ZN(n_0_0_132));
   AOI21_X1 i_0_0_297 (.A(n_0_0_134), .B1(n_0_0_136), .B2(n_0_0_135), .ZN(
      n_0_0_133));
   NOR2_X1 i_0_0_298 (.A1(n_0_0_206), .A2(end_T_address[15]), .ZN(n_0_0_134));
   AOI22_X1 i_0_0_299 (.A1(end_T_address[15]), .A2(n_0_0_206), .B1(n_0_0_205), 
      .B2(end_T_address[14]), .ZN(n_0_0_135));
   OAI221_X1 i_0_0_300 (.A(n_0_0_137), .B1(n_0_0_204), .B2(end_T_address[13]), 
      .C1(end_T_address[14]), .C2(n_0_0_205), .ZN(n_0_0_136));
   NAND2_X1 i_0_0_301 (.A1(n_0_0_139), .A2(n_0_0_138), .ZN(n_0_0_137));
   AOI22_X1 i_0_0_302 (.A1(end_T_address[13]), .A2(n_0_0_204), .B1(n_0_0_203), 
      .B2(end_T_address[12]), .ZN(n_0_0_138));
   OAI21_X1 i_0_0_303 (.A(n_0_0_140), .B1(n_0_0_203), .B2(end_T_address[12]), 
      .ZN(n_0_0_139));
   AOI21_X1 i_0_0_304 (.A(n_0_0_141), .B1(n_0_0_143), .B2(n_0_0_142), .ZN(
      n_0_0_140));
   NOR2_X1 i_0_0_305 (.A1(n_0_0_202), .A2(end_T_address[11]), .ZN(n_0_0_141));
   AOI22_X1 i_0_0_306 (.A1(end_T_address[11]), .A2(n_0_0_202), .B1(n_0_0_201), 
      .B2(end_T_address[10]), .ZN(n_0_0_142));
   OAI221_X1 i_0_0_307 (.A(n_0_0_144), .B1(n_0_0_200), .B2(end_T_address[9]), 
      .C1(end_T_address[10]), .C2(n_0_0_201), .ZN(n_0_0_143));
   NAND2_X1 i_0_0_308 (.A1(n_0_0_146), .A2(n_0_0_145), .ZN(n_0_0_144));
   AOI22_X1 i_0_0_309 (.A1(end_T_address[9]), .A2(n_0_0_200), .B1(n_0_0_199), 
      .B2(end_T_address[8]), .ZN(n_0_0_145));
   OAI21_X1 i_0_0_310 (.A(n_0_0_147), .B1(n_0_0_199), .B2(end_T_address[8]), 
      .ZN(n_0_0_146));
   AOI21_X1 i_0_0_311 (.A(n_0_0_148), .B1(n_0_0_150), .B2(n_0_0_149), .ZN(
      n_0_0_147));
   NOR2_X1 i_0_0_312 (.A1(n_0_0_198), .A2(end_T_address[7]), .ZN(n_0_0_148));
   AOI22_X1 i_0_0_313 (.A1(end_T_address[7]), .A2(n_0_0_198), .B1(n_0_0_197), 
      .B2(end_T_address[6]), .ZN(n_0_0_149));
   OAI221_X1 i_0_0_314 (.A(n_0_0_151), .B1(n_0_0_196), .B2(end_T_address[5]), 
      .C1(end_T_address[6]), .C2(n_0_0_197), .ZN(n_0_0_150));
   OAI21_X1 i_0_0_315 (.A(n_0_0_152), .B1(n_0_0_154), .B2(n_0_0_153), .ZN(
      n_0_0_151));
   AOI22_X1 i_0_0_316 (.A1(end_T_address[5]), .A2(n_0_0_196), .B1(n_0_0_195), 
      .B2(end_T_address[4]), .ZN(n_0_0_152));
   OAI22_X1 i_0_0_317 (.A1(end_T_address[4]), .A2(n_0_0_195), .B1(n_0_0_194), 
      .B2(end_T_address[3]), .ZN(n_0_0_153));
   AOI221_X1 i_0_0_318 (.A(n_0_0_155), .B1(n_0_0_193), .B2(end_T_address[2]), 
      .C1(end_T_address[3]), .C2(n_0_0_194), .ZN(n_0_0_154));
   NOR2_X1 i_0_0_319 (.A1(n_0_0_157), .A2(n_0_0_156), .ZN(n_0_0_155));
   OAI22_X1 i_0_0_320 (.A1(end_T_address[2]), .A2(n_0_0_193), .B1(n_0_0_192), 
      .B2(end_T_address[1]), .ZN(n_0_0_156));
   AOI22_X1 i_0_0_321 (.A1(end_T_address[1]), .A2(n_0_0_192), .B1(n_0_0_191), 
      .B2(end_T_address[0]), .ZN(n_0_0_157));
   NOR2_X1 i_0_0_322 (.A1(enable_output_IO), .A2(RST), .ZN(n_0_295));
   INV_X1 i_0_0_323 (.A(CLK), .ZN(n_0_201));
   INV_X1 i_0_0_324 (.A(state_reg[1]), .ZN(n_0_0_158));
   INV_X1 i_0_0_325 (.A(RST), .ZN(n_0_0_159));
   INV_X1 i_0_0_326 (.A(n_0_47), .ZN(n_0_0_160));
   INV_X1 i_0_0_327 (.A(n_0_46), .ZN(n_0_0_161));
   INV_X1 i_0_0_328 (.A(n_0_43), .ZN(n_0_0_162));
   INV_X1 i_0_0_329 (.A(n_0_42), .ZN(n_0_0_163));
   INV_X1 i_0_0_330 (.A(n_0_39), .ZN(n_0_0_164));
   INV_X1 i_0_0_331 (.A(n_0_38), .ZN(n_0_0_165));
   INV_X1 i_0_0_332 (.A(n_0_2), .ZN(n_0_0_166));
   INV_X1 i_0_0_333 (.A(n_0_1), .ZN(n_0_0_167));
   INV_X1 i_0_0_334 (.A(n_0_292), .ZN(n_0_0_168));
   INV_X1 i_0_0_335 (.A(n_0_290), .ZN(n_0_0_169));
   INV_X1 i_0_0_336 (.A(n_0_284), .ZN(n_0_0_170));
   INV_X1 i_0_0_337 (.A(n_0_282), .ZN(n_0_0_171));
   INV_X1 i_0_0_338 (.A(n_0_276), .ZN(n_0_0_172));
   INV_X1 i_0_0_339 (.A(n_0_274), .ZN(n_0_0_173));
   INV_X1 i_0_0_340 (.A(n_0_272), .ZN(n_0_0_174));
   INV_X1 i_0_0_341 (.A(end_Output_address[1]), .ZN(n_0_0_175));
   INV_X1 i_0_0_342 (.A(end_Output_address[2]), .ZN(n_0_0_176));
   INV_X1 i_0_0_343 (.A(end_Output_address[3]), .ZN(n_0_0_177));
   INV_X1 i_0_0_344 (.A(end_Output_address[6]), .ZN(n_0_0_178));
   INV_X1 i_0_0_345 (.A(end_Output_address[7]), .ZN(n_0_0_179));
   INV_X1 i_0_0_346 (.A(end_Output_address[10]), .ZN(n_0_0_180));
   INV_X1 i_0_0_347 (.A(end_Output_address[11]), .ZN(n_0_0_181));
   INV_X1 i_0_0_348 (.A(end_Output_address[14]), .ZN(n_0_0_182));
   INV_X1 i_0_0_349 (.A(end_Output_address[15]), .ZN(n_0_0_183));
   INV_X1 i_0_0_350 (.A(end_Output_address[18]), .ZN(n_0_0_184));
   INV_X1 i_0_0_351 (.A(end_Output_address[19]), .ZN(n_0_0_185));
   INV_X1 i_0_0_352 (.A(end_Output_address[22]), .ZN(n_0_0_186));
   INV_X1 i_0_0_353 (.A(end_Output_address[23]), .ZN(n_0_0_187));
   INV_X1 i_0_0_354 (.A(end_Output_address[26]), .ZN(n_0_0_188));
   INV_X1 i_0_0_355 (.A(end_Output_address[27]), .ZN(n_0_0_189));
   INV_X1 i_0_0_356 (.A(end_Output_address[31]), .ZN(n_0_0_190));
   INV_X1 i_0_0_357 (.A(n_0_116), .ZN(n_0_0_191));
   INV_X1 i_0_0_358 (.A(n_0_115), .ZN(n_0_0_192));
   INV_X1 i_0_0_359 (.A(n_0_114), .ZN(n_0_0_193));
   INV_X1 i_0_0_360 (.A(n_0_113), .ZN(n_0_0_194));
   INV_X1 i_0_0_361 (.A(n_0_112), .ZN(n_0_0_195));
   INV_X1 i_0_0_362 (.A(n_0_111), .ZN(n_0_0_196));
   INV_X1 i_0_0_363 (.A(n_0_110), .ZN(n_0_0_197));
   INV_X1 i_0_0_364 (.A(n_0_109), .ZN(n_0_0_198));
   INV_X1 i_0_0_365 (.A(n_0_108), .ZN(n_0_0_199));
   INV_X1 i_0_0_366 (.A(n_0_107), .ZN(n_0_0_200));
   INV_X1 i_0_0_367 (.A(n_0_106), .ZN(n_0_0_201));
   INV_X1 i_0_0_368 (.A(n_0_105), .ZN(n_0_0_202));
   INV_X1 i_0_0_369 (.A(n_0_104), .ZN(n_0_0_203));
   INV_X1 i_0_0_370 (.A(n_0_103), .ZN(n_0_0_204));
   INV_X1 i_0_0_371 (.A(n_0_102), .ZN(n_0_0_205));
   INV_X1 i_0_0_372 (.A(n_0_101), .ZN(n_0_0_206));
   INV_X1 i_0_0_373 (.A(n_0_100), .ZN(n_0_0_207));
   INV_X1 i_0_0_374 (.A(n_0_99), .ZN(n_0_0_208));
   INV_X1 i_0_0_375 (.A(n_0_98), .ZN(n_0_0_209));
   INV_X1 i_0_0_376 (.A(n_0_97), .ZN(n_0_0_210));
   INV_X1 i_0_0_377 (.A(n_0_96), .ZN(n_0_0_211));
   INV_X1 i_0_0_378 (.A(n_0_95), .ZN(n_0_0_212));
   INV_X1 i_0_0_379 (.A(n_0_94), .ZN(n_0_0_213));
   INV_X1 i_0_0_380 (.A(n_0_93), .ZN(n_0_0_214));
   INV_X1 i_0_0_381 (.A(n_0_92), .ZN(n_0_0_215));
   INV_X1 i_0_0_382 (.A(n_0_91), .ZN(n_0_0_216));
   INV_X1 i_0_0_383 (.A(n_0_90), .ZN(n_0_0_217));
   INV_X1 i_0_0_384 (.A(n_0_89), .ZN(n_0_0_218));
   INV_X1 i_0_0_385 (.A(n_0_88), .ZN(n_0_0_219));
   INV_X1 i_0_0_386 (.A(n_0_87), .ZN(n_0_0_220));
   INV_X1 i_0_0_387 (.A(n_0_86), .ZN(n_0_0_221));
   INV_X1 i_0_0_388 (.A(end_T_address[31]), .ZN(n_0_0_222));
endmodule
